magic
tech scmos
timestamp 1619104829
<< nwell >>
rect 143 1875 169 1901
rect 233 1875 259 1901
rect 42 1803 68 1829
rect 143 1823 169 1849
rect 233 1823 259 1849
rect 77 1792 103 1818
rect -176 1739 -150 1765
rect -137 1739 -111 1765
rect -97 1739 -71 1765
rect -58 1739 -32 1765
rect -17 1739 9 1765
rect 42 1751 68 1777
rect 147 1745 173 1771
rect 237 1745 263 1771
rect -188 1681 -162 1707
rect 147 1693 173 1719
rect 237 1693 263 1719
rect 143 1619 169 1645
rect 233 1619 259 1645
rect 42 1547 68 1573
rect 143 1567 169 1593
rect 233 1567 259 1593
rect 77 1536 103 1562
rect -176 1483 -150 1509
rect -137 1483 -111 1509
rect -97 1483 -71 1509
rect -58 1483 -32 1509
rect -17 1483 9 1509
rect 42 1495 68 1521
rect 147 1489 173 1515
rect 237 1489 263 1515
rect 313 1512 339 1538
rect 1325 1520 1351 1546
rect 1415 1520 1441 1546
rect 399 1482 425 1508
rect -188 1425 -162 1451
rect 147 1437 173 1463
rect 237 1437 263 1463
rect 339 1410 365 1436
rect 399 1430 425 1456
rect 485 1437 511 1463
rect 1224 1448 1250 1474
rect 1325 1468 1351 1494
rect 1415 1468 1441 1494
rect 1259 1437 1285 1463
rect 143 1363 169 1389
rect 233 1363 259 1389
rect 399 1387 425 1413
rect 485 1385 511 1411
rect 773 1370 799 1396
rect 1006 1384 1032 1410
rect 1045 1384 1071 1410
rect 1085 1384 1111 1410
rect 1124 1384 1150 1410
rect 1165 1384 1191 1410
rect 1224 1396 1250 1422
rect 1329 1390 1355 1416
rect 1419 1390 1445 1416
rect 42 1291 68 1317
rect 143 1311 169 1337
rect 233 1311 259 1337
rect 399 1335 425 1361
rect 859 1340 885 1366
rect 994 1326 1020 1352
rect 1329 1338 1355 1364
rect 1419 1338 1445 1364
rect 77 1280 103 1306
rect 354 1274 380 1300
rect 390 1266 416 1292
rect 799 1268 825 1294
rect 859 1288 885 1314
rect 945 1295 971 1321
rect -176 1227 -150 1253
rect -137 1227 -111 1253
rect -97 1227 -71 1253
rect -58 1227 -32 1253
rect -17 1227 9 1253
rect 42 1239 68 1265
rect 147 1233 173 1259
rect 237 1233 263 1259
rect 354 1222 380 1248
rect 859 1245 885 1271
rect 945 1243 971 1269
rect 1325 1264 1351 1290
rect 1415 1264 1441 1290
rect -188 1169 -162 1195
rect 147 1181 173 1207
rect 237 1181 263 1207
rect 313 1177 339 1203
rect 859 1193 885 1219
rect 1224 1192 1250 1218
rect 1325 1212 1351 1238
rect 1415 1212 1441 1238
rect 1259 1181 1285 1207
rect 399 1147 425 1173
rect 773 1137 799 1163
rect 143 1107 169 1133
rect 233 1107 259 1133
rect 42 1035 68 1061
rect 143 1055 169 1081
rect 233 1055 259 1081
rect 339 1075 365 1101
rect 399 1095 425 1121
rect 485 1102 511 1128
rect 859 1107 885 1133
rect 1006 1128 1032 1154
rect 1045 1128 1071 1154
rect 1085 1128 1111 1154
rect 1124 1128 1150 1154
rect 1165 1128 1191 1154
rect 1224 1140 1250 1166
rect 1329 1134 1355 1160
rect 1419 1134 1445 1160
rect 399 1052 425 1078
rect 485 1050 511 1076
rect 77 1024 103 1050
rect -176 971 -150 997
rect -137 971 -111 997
rect -97 971 -71 997
rect -58 971 -32 997
rect -17 971 9 997
rect 42 983 68 1009
rect 147 977 173 1003
rect 237 977 263 1003
rect 399 1000 425 1026
rect 535 1017 561 1043
rect 573 1017 599 1043
rect 611 1017 637 1043
rect 649 1017 675 1043
rect 718 1018 744 1044
rect 799 1035 825 1061
rect 859 1055 885 1081
rect 945 1062 971 1088
rect 994 1070 1020 1096
rect 1329 1082 1355 1108
rect 1419 1082 1445 1108
rect 859 1012 885 1038
rect 945 1010 971 1036
rect 1325 1008 1351 1034
rect 1415 1008 1441 1034
rect -188 913 -162 939
rect 147 925 173 951
rect 237 925 263 951
rect 354 939 380 965
rect 718 961 744 987
rect 859 960 885 986
rect 390 931 416 957
rect 1224 936 1250 962
rect 1325 956 1351 982
rect 1415 956 1441 982
rect 354 887 380 913
rect 718 904 744 930
rect 773 904 799 930
rect 1259 925 1285 951
rect 143 851 169 877
rect 233 851 259 877
rect 859 874 885 900
rect 313 842 339 868
rect 718 847 744 873
rect 1006 872 1032 898
rect 1045 872 1071 898
rect 1085 872 1111 898
rect 1124 872 1150 898
rect 1165 872 1191 898
rect 1224 884 1250 910
rect 1329 878 1355 904
rect 1419 878 1445 904
rect 42 779 68 805
rect 143 799 169 825
rect 233 799 259 825
rect 399 812 425 838
rect 799 802 825 828
rect 859 822 885 848
rect 945 829 971 855
rect 994 814 1020 840
rect 1329 826 1355 852
rect 1419 826 1445 852
rect 77 768 103 794
rect -176 715 -150 741
rect -137 715 -111 741
rect -97 715 -71 741
rect -58 715 -32 741
rect -17 715 9 741
rect 42 727 68 753
rect 147 721 173 747
rect 237 721 263 747
rect 339 740 365 766
rect 399 760 425 786
rect 485 767 511 793
rect 859 779 885 805
rect 945 777 971 803
rect 399 717 425 743
rect 485 715 511 741
rect 859 727 885 753
rect 1325 752 1351 778
rect 1415 752 1441 778
rect -188 657 -162 683
rect 147 669 173 695
rect 237 669 263 695
rect 399 665 425 691
rect 773 671 799 697
rect 1224 680 1250 706
rect 1325 700 1351 726
rect 1415 700 1441 726
rect 1259 669 1285 695
rect 859 641 885 667
rect 143 595 169 621
rect 233 595 259 621
rect 354 604 380 630
rect 390 596 416 622
rect 42 523 68 549
rect 143 543 169 569
rect 233 543 259 569
rect 354 552 380 578
rect 799 569 825 595
rect 859 589 885 615
rect 945 596 971 622
rect 1006 616 1032 642
rect 1045 616 1071 642
rect 1085 616 1111 642
rect 1124 616 1150 642
rect 1165 616 1191 642
rect 1224 628 1250 654
rect 1329 622 1355 648
rect 1419 622 1445 648
rect 859 546 885 572
rect 945 544 971 570
rect 994 558 1020 584
rect 1329 570 1355 596
rect 1419 570 1445 596
rect 77 512 103 538
rect 313 507 339 533
rect -176 459 -150 485
rect -137 459 -111 485
rect -97 459 -71 485
rect -58 459 -32 485
rect -17 459 9 485
rect 42 471 68 497
rect 147 465 173 491
rect 237 465 263 491
rect 399 477 425 503
rect 773 495 799 521
rect 859 494 885 520
rect 1325 496 1351 522
rect 1415 496 1441 522
rect -188 401 -162 427
rect 147 413 173 439
rect 237 413 263 439
rect 339 405 365 431
rect 399 425 425 451
rect 485 432 511 458
rect 1224 424 1250 450
rect 1325 444 1351 470
rect 1415 444 1441 470
rect 1259 413 1285 439
rect 399 382 425 408
rect 485 380 511 406
rect 143 339 169 365
rect 233 339 259 365
rect 1006 360 1032 386
rect 1045 360 1071 386
rect 1085 360 1111 386
rect 1124 360 1150 386
rect 1165 360 1191 386
rect 1224 372 1250 398
rect 1329 366 1355 392
rect 1419 366 1445 392
rect 399 330 425 356
rect 42 267 68 293
rect 143 287 169 313
rect 233 287 259 313
rect 994 302 1020 328
rect 1329 314 1355 340
rect 1419 314 1445 340
rect 77 256 103 282
rect 354 269 380 295
rect 390 261 416 287
rect -176 203 -150 229
rect -137 203 -111 229
rect -97 203 -71 229
rect -58 203 -32 229
rect -17 203 9 229
rect 42 215 68 241
rect 147 209 173 235
rect 237 209 263 235
rect 354 217 380 243
rect -188 145 -162 171
rect 147 157 173 183
rect 237 157 263 183
rect 143 83 169 109
rect 233 83 259 109
rect 42 11 68 37
rect 143 31 169 57
rect 233 31 259 57
rect 77 0 103 26
rect -176 -53 -150 -27
rect -137 -53 -111 -27
rect -97 -53 -71 -27
rect -58 -53 -32 -27
rect -17 -53 9 -27
rect 42 -41 68 -15
rect 147 -47 173 -21
rect 237 -47 263 -21
rect -188 -111 -162 -85
rect 147 -99 173 -73
rect 237 -99 263 -73
<< ntransistor >>
rect 103 1869 111 1871
rect 193 1869 201 1871
rect 125 1861 133 1863
rect 215 1861 223 1863
rect 2 1797 10 1799
rect 24 1789 32 1791
rect 89 1778 91 1786
rect 107 1739 115 1741
rect 197 1739 205 1741
rect -164 1725 -162 1733
rect -125 1725 -123 1733
rect -85 1725 -83 1733
rect -46 1725 -44 1733
rect -5 1725 -3 1733
rect 129 1731 137 1733
rect 219 1731 227 1733
rect -176 1667 -174 1675
rect 103 1613 111 1615
rect 193 1613 201 1615
rect 125 1605 133 1607
rect 215 1605 223 1607
rect 2 1541 10 1543
rect 24 1533 32 1535
rect 89 1522 91 1530
rect 1285 1514 1293 1516
rect 1375 1514 1383 1516
rect 1307 1506 1315 1508
rect 1397 1506 1405 1508
rect 325 1498 327 1506
rect 107 1483 115 1485
rect 197 1483 205 1485
rect -164 1469 -162 1477
rect -125 1469 -123 1477
rect -85 1469 -83 1477
rect -46 1469 -44 1477
rect -5 1469 -3 1477
rect 129 1475 137 1477
rect 219 1475 227 1477
rect 359 1476 367 1478
rect 381 1468 389 1470
rect 1184 1442 1192 1444
rect 1206 1434 1214 1436
rect 445 1431 453 1433
rect 325 1422 333 1424
rect 467 1423 475 1425
rect -176 1411 -174 1419
rect 1271 1423 1273 1431
rect 359 1381 367 1383
rect 1289 1384 1297 1386
rect 1379 1384 1387 1386
rect 381 1373 389 1375
rect 1018 1370 1020 1378
rect 1057 1370 1059 1378
rect 1097 1370 1099 1378
rect 1136 1370 1138 1378
rect 1177 1370 1179 1378
rect 1311 1376 1319 1378
rect 1401 1376 1409 1378
rect 103 1357 111 1359
rect 193 1357 201 1359
rect 785 1356 787 1364
rect 125 1349 133 1351
rect 215 1349 223 1351
rect 819 1334 827 1336
rect 841 1326 849 1328
rect 1006 1312 1008 1320
rect 2 1285 10 1287
rect 24 1277 32 1279
rect 905 1289 913 1291
rect 785 1280 793 1282
rect 927 1281 935 1283
rect 89 1266 91 1274
rect 314 1268 322 1270
rect 336 1260 344 1262
rect 402 1252 404 1260
rect 1285 1258 1293 1260
rect 1375 1258 1383 1260
rect 1307 1250 1315 1252
rect 1397 1250 1405 1252
rect 819 1239 827 1241
rect 107 1227 115 1229
rect 197 1227 205 1229
rect 841 1231 849 1233
rect -164 1213 -162 1221
rect -125 1213 -123 1221
rect -85 1213 -83 1221
rect -46 1213 -44 1221
rect -5 1213 -3 1221
rect 129 1219 137 1221
rect 219 1219 227 1221
rect 1184 1186 1192 1188
rect 1206 1178 1214 1180
rect 325 1163 327 1171
rect -176 1155 -174 1163
rect 1271 1167 1273 1175
rect 359 1141 367 1143
rect 381 1133 389 1135
rect 785 1123 787 1131
rect 1289 1128 1297 1130
rect 1379 1128 1387 1130
rect 1018 1114 1020 1122
rect 1057 1114 1059 1122
rect 1097 1114 1099 1122
rect 1136 1114 1138 1122
rect 1177 1114 1179 1122
rect 1311 1120 1319 1122
rect 1401 1120 1409 1122
rect 103 1101 111 1103
rect 193 1101 201 1103
rect 819 1101 827 1103
rect 125 1093 133 1095
rect 215 1093 223 1095
rect 445 1096 453 1098
rect 841 1093 849 1095
rect 325 1087 333 1089
rect 467 1088 475 1090
rect 905 1056 913 1058
rect 1006 1056 1008 1064
rect 359 1046 367 1048
rect 785 1047 793 1049
rect 927 1048 935 1050
rect 381 1038 389 1040
rect 2 1029 10 1031
rect 24 1021 32 1023
rect 89 1010 91 1018
rect 730 1004 732 1012
rect 819 1006 827 1008
rect 1285 1002 1293 1004
rect 1375 1002 1383 1004
rect 841 998 849 1000
rect 661 983 663 991
rect 691 984 693 992
rect 1307 994 1315 996
rect 1397 994 1405 996
rect 107 971 115 973
rect 197 971 205 973
rect -164 957 -162 965
rect -125 957 -123 965
rect -85 957 -83 965
rect -46 957 -44 965
rect -5 957 -3 965
rect 129 963 137 965
rect 219 963 227 965
rect 653 953 655 961
rect 623 942 625 950
rect 730 947 732 955
rect 314 933 322 935
rect 336 925 344 927
rect 1184 930 1192 932
rect 402 917 404 925
rect 1206 922 1214 924
rect 615 912 617 920
rect -176 899 -174 907
rect 585 901 587 909
rect 1271 911 1273 919
rect 730 890 732 898
rect 785 890 787 898
rect 577 871 579 879
rect 819 868 827 870
rect 547 860 549 868
rect 1289 872 1297 874
rect 1379 872 1387 874
rect 841 860 849 862
rect 103 845 111 847
rect 193 845 201 847
rect 125 837 133 839
rect 215 837 223 839
rect 1018 858 1020 866
rect 1057 858 1059 866
rect 1097 858 1099 866
rect 1136 858 1138 866
rect 1177 858 1179 866
rect 1311 864 1319 866
rect 1401 864 1409 866
rect 325 828 327 836
rect 539 831 541 839
rect 730 833 732 841
rect 905 823 913 825
rect 785 814 793 816
rect 927 815 935 817
rect 359 806 367 808
rect 531 802 533 810
rect 381 798 389 800
rect 1006 800 1008 808
rect 2 773 10 775
rect 24 765 32 767
rect 819 773 827 775
rect 841 765 849 767
rect 89 754 91 762
rect 445 761 453 763
rect 325 752 333 754
rect 467 753 475 755
rect 1285 746 1293 748
rect 1375 746 1383 748
rect 1307 738 1315 740
rect 1397 738 1405 740
rect 107 715 115 717
rect 197 715 205 717
rect 359 711 367 713
rect -164 701 -162 709
rect -125 701 -123 709
rect -85 701 -83 709
rect -46 701 -44 709
rect -5 701 -3 709
rect 129 707 137 709
rect 219 707 227 709
rect 381 703 389 705
rect 1184 674 1192 676
rect 1206 666 1214 668
rect 785 657 787 665
rect 1271 655 1273 663
rect -176 643 -174 651
rect 819 635 827 637
rect 841 627 849 629
rect 1289 616 1297 618
rect 1379 616 1387 618
rect 314 598 322 600
rect 103 589 111 591
rect 193 589 201 591
rect 336 590 344 592
rect 1018 602 1020 610
rect 1057 602 1059 610
rect 1097 602 1099 610
rect 1136 602 1138 610
rect 1177 602 1179 610
rect 1311 608 1319 610
rect 1401 608 1409 610
rect 125 581 133 583
rect 215 581 223 583
rect 402 582 404 590
rect 905 590 913 592
rect 785 581 793 583
rect 927 582 935 584
rect 1006 544 1008 552
rect 819 540 827 542
rect 841 532 849 534
rect 2 517 10 519
rect 24 509 32 511
rect 89 498 91 506
rect 325 493 327 501
rect 1285 490 1293 492
rect 1375 490 1383 492
rect 785 481 787 489
rect 1307 482 1315 484
rect 1397 482 1405 484
rect 359 471 367 473
rect 381 463 389 465
rect 107 459 115 461
rect 197 459 205 461
rect -164 445 -162 453
rect -125 445 -123 453
rect -85 445 -83 453
rect -46 445 -44 453
rect -5 445 -3 453
rect 129 451 137 453
rect 219 451 227 453
rect 445 426 453 428
rect 325 417 333 419
rect 467 418 475 420
rect 1184 418 1192 420
rect 1206 410 1214 412
rect -176 387 -174 395
rect 1271 399 1273 407
rect 359 376 367 378
rect 381 368 389 370
rect 1289 360 1297 362
rect 1379 360 1387 362
rect 1018 346 1020 354
rect 1057 346 1059 354
rect 1097 346 1099 354
rect 1136 346 1138 354
rect 1177 346 1179 354
rect 1311 352 1319 354
rect 1401 352 1409 354
rect 103 333 111 335
rect 193 333 201 335
rect 125 325 133 327
rect 215 325 223 327
rect 1006 288 1008 296
rect 2 261 10 263
rect 314 263 322 265
rect 24 253 32 255
rect 336 255 344 257
rect 89 242 91 250
rect 402 247 404 255
rect 107 203 115 205
rect 197 203 205 205
rect -164 189 -162 197
rect -125 189 -123 197
rect -85 189 -83 197
rect -46 189 -44 197
rect -5 189 -3 197
rect 129 195 137 197
rect 219 195 227 197
rect -176 131 -174 139
rect 103 77 111 79
rect 193 77 201 79
rect 125 69 133 71
rect 215 69 223 71
rect 2 5 10 7
rect 24 -3 32 -1
rect 89 -14 91 -6
rect 107 -53 115 -51
rect 197 -53 205 -51
rect -164 -67 -162 -59
rect -125 -67 -123 -59
rect -85 -67 -83 -59
rect -46 -67 -44 -59
rect -5 -67 -3 -59
rect 129 -61 137 -59
rect 219 -61 227 -59
rect -176 -125 -174 -117
<< ptransistor >>
rect 149 1887 157 1889
rect 239 1887 247 1889
rect 149 1835 157 1837
rect 239 1835 247 1837
rect 48 1815 56 1817
rect 89 1798 91 1806
rect 48 1763 56 1765
rect 153 1757 161 1759
rect 243 1757 251 1759
rect -164 1745 -162 1753
rect -125 1745 -123 1753
rect -85 1745 -83 1753
rect -46 1745 -44 1753
rect -5 1745 -3 1753
rect 153 1705 161 1707
rect 243 1705 251 1707
rect -176 1687 -174 1695
rect 149 1631 157 1633
rect 239 1631 247 1633
rect 149 1579 157 1581
rect 239 1579 247 1581
rect 48 1559 56 1561
rect 89 1542 91 1550
rect 1331 1532 1339 1534
rect 1421 1532 1429 1534
rect 325 1518 327 1526
rect 48 1507 56 1509
rect 153 1501 161 1503
rect 243 1501 251 1503
rect -164 1489 -162 1497
rect -125 1489 -123 1497
rect -85 1489 -83 1497
rect -46 1489 -44 1497
rect -5 1489 -3 1497
rect 405 1494 413 1496
rect 1331 1480 1339 1482
rect 1421 1480 1429 1482
rect 1230 1460 1238 1462
rect 153 1449 161 1451
rect 243 1449 251 1451
rect 491 1449 499 1451
rect 405 1442 413 1444
rect -176 1431 -174 1439
rect 1271 1443 1273 1451
rect 345 1422 353 1424
rect 1230 1408 1238 1410
rect 405 1399 413 1401
rect 491 1397 499 1399
rect 1335 1402 1343 1404
rect 1425 1402 1433 1404
rect 1018 1390 1020 1398
rect 1057 1390 1059 1398
rect 1097 1390 1099 1398
rect 1136 1390 1138 1398
rect 1177 1390 1179 1398
rect 149 1375 157 1377
rect 239 1375 247 1377
rect 785 1376 787 1384
rect 865 1352 873 1354
rect 405 1347 413 1349
rect 1335 1350 1343 1352
rect 1425 1350 1433 1352
rect 1006 1332 1008 1340
rect 149 1323 157 1325
rect 239 1323 247 1325
rect 951 1307 959 1309
rect 48 1303 56 1305
rect 865 1300 873 1302
rect 89 1286 91 1294
rect 360 1286 368 1288
rect 805 1280 813 1282
rect 402 1272 404 1280
rect 1331 1276 1339 1278
rect 1421 1276 1429 1278
rect 48 1251 56 1253
rect 865 1257 873 1259
rect 951 1255 959 1257
rect 153 1245 161 1247
rect 243 1245 251 1247
rect -164 1233 -162 1241
rect -125 1233 -123 1241
rect -85 1233 -83 1241
rect -46 1233 -44 1241
rect -5 1233 -3 1241
rect 360 1234 368 1236
rect 1331 1224 1339 1226
rect 1421 1224 1429 1226
rect 865 1205 873 1207
rect 1230 1204 1238 1206
rect 153 1193 161 1195
rect 243 1193 251 1195
rect 325 1183 327 1191
rect 1271 1187 1273 1195
rect -176 1175 -174 1183
rect 405 1159 413 1161
rect 1230 1152 1238 1154
rect 785 1143 787 1151
rect 1335 1146 1343 1148
rect 1425 1146 1433 1148
rect 1018 1134 1020 1142
rect 1057 1134 1059 1142
rect 1097 1134 1099 1142
rect 1136 1134 1138 1142
rect 1177 1134 1179 1142
rect 149 1119 157 1121
rect 239 1119 247 1121
rect 865 1119 873 1121
rect 491 1114 499 1116
rect 405 1107 413 1109
rect 1335 1094 1343 1096
rect 1425 1094 1433 1096
rect 345 1087 353 1089
rect 1006 1076 1008 1084
rect 951 1074 959 1076
rect 149 1067 157 1069
rect 239 1067 247 1069
rect 405 1064 413 1066
rect 865 1067 873 1069
rect 491 1062 499 1064
rect 48 1047 56 1049
rect 805 1047 813 1049
rect 89 1030 91 1038
rect 547 1023 549 1031
rect 585 1023 587 1031
rect 623 1023 625 1031
rect 661 1023 663 1031
rect 730 1024 732 1032
rect 865 1024 873 1026
rect 405 1012 413 1014
rect 951 1022 959 1024
rect 1331 1020 1339 1022
rect 1421 1020 1429 1022
rect 48 995 56 997
rect 153 989 161 991
rect 243 989 251 991
rect -164 977 -162 985
rect -125 977 -123 985
rect -85 977 -83 985
rect -46 977 -44 985
rect -5 977 -3 985
rect 730 967 732 975
rect 865 972 873 974
rect 1331 968 1339 970
rect 1421 968 1429 970
rect 360 951 368 953
rect 153 937 161 939
rect 243 937 251 939
rect 402 937 404 945
rect 1230 948 1238 950
rect -176 919 -174 927
rect 1271 931 1273 939
rect 730 910 732 918
rect 785 910 787 918
rect 360 899 368 901
rect 1230 896 1238 898
rect 865 886 873 888
rect 1335 890 1343 892
rect 1425 890 1433 892
rect 1018 878 1020 886
rect 1057 878 1059 886
rect 1097 878 1099 886
rect 1136 878 1138 886
rect 1177 878 1179 886
rect 149 863 157 865
rect 239 863 247 865
rect 325 848 327 856
rect 730 853 732 861
rect 951 841 959 843
rect 1335 838 1343 840
rect 1425 838 1433 840
rect 865 834 873 836
rect 405 824 413 826
rect 1006 820 1008 828
rect 149 811 157 813
rect 239 811 247 813
rect 805 814 813 816
rect 48 791 56 793
rect 865 791 873 793
rect 951 789 959 791
rect 89 774 91 782
rect 491 779 499 781
rect 405 772 413 774
rect 1331 764 1339 766
rect 1421 764 1429 766
rect 345 752 353 754
rect 48 739 56 741
rect 865 739 873 741
rect 153 733 161 735
rect 243 733 251 735
rect -164 721 -162 729
rect -125 721 -123 729
rect -85 721 -83 729
rect -46 721 -44 729
rect -5 721 -3 729
rect 405 729 413 731
rect 491 727 499 729
rect 1331 712 1339 714
rect 1421 712 1429 714
rect 1230 692 1238 694
rect 153 681 161 683
rect 243 681 251 683
rect 405 677 413 679
rect 785 677 787 685
rect -176 663 -174 671
rect 1271 675 1273 683
rect 865 653 873 655
rect 1230 640 1238 642
rect 1335 634 1343 636
rect 1425 634 1433 636
rect 1018 622 1020 630
rect 1057 622 1059 630
rect 1097 622 1099 630
rect 1136 622 1138 630
rect 1177 622 1179 630
rect 360 616 368 618
rect 149 607 157 609
rect 239 607 247 609
rect 402 602 404 610
rect 951 608 959 610
rect 865 601 873 603
rect 805 581 813 583
rect 1335 582 1343 584
rect 1425 582 1433 584
rect 360 564 368 566
rect 149 555 157 557
rect 239 555 247 557
rect 1006 564 1008 572
rect 865 558 873 560
rect 951 556 959 558
rect 48 535 56 537
rect 89 518 91 526
rect 325 513 327 521
rect 785 501 787 509
rect 1331 508 1339 510
rect 1421 508 1429 510
rect 865 506 873 508
rect 405 489 413 491
rect 48 483 56 485
rect 153 477 161 479
rect 243 477 251 479
rect -164 465 -162 473
rect -125 465 -123 473
rect -85 465 -83 473
rect -46 465 -44 473
rect -5 465 -3 473
rect 1331 456 1339 458
rect 1421 456 1429 458
rect 491 444 499 446
rect 405 437 413 439
rect 1230 436 1238 438
rect 153 425 161 427
rect 243 425 251 427
rect 345 417 353 419
rect 1271 419 1273 427
rect -176 407 -174 415
rect 405 394 413 396
rect 491 392 499 394
rect 1230 384 1238 386
rect 1335 378 1343 380
rect 1425 378 1433 380
rect 1018 366 1020 374
rect 1057 366 1059 374
rect 1097 366 1099 374
rect 1136 366 1138 374
rect 1177 366 1179 374
rect 149 351 157 353
rect 239 351 247 353
rect 405 342 413 344
rect 1335 326 1343 328
rect 1425 326 1433 328
rect 1006 308 1008 316
rect 149 299 157 301
rect 239 299 247 301
rect 360 281 368 283
rect 48 279 56 281
rect 89 262 91 270
rect 402 267 404 275
rect 48 227 56 229
rect 360 229 368 231
rect 153 221 161 223
rect 243 221 251 223
rect -164 209 -162 217
rect -125 209 -123 217
rect -85 209 -83 217
rect -46 209 -44 217
rect -5 209 -3 217
rect 153 169 161 171
rect 243 169 251 171
rect -176 151 -174 159
rect 149 95 157 97
rect 239 95 247 97
rect 149 43 157 45
rect 239 43 247 45
rect 48 23 56 25
rect 89 6 91 14
rect 48 -29 56 -27
rect 153 -35 161 -33
rect 243 -35 251 -33
rect -164 -47 -162 -39
rect -125 -47 -123 -39
rect -85 -47 -83 -39
rect -46 -47 -44 -39
rect -5 -47 -3 -39
rect 153 -87 161 -85
rect 243 -87 251 -85
rect -176 -105 -174 -97
<< ndiffusion >>
rect 103 1871 111 1872
rect 193 1871 201 1872
rect 103 1868 111 1869
rect 193 1868 201 1869
rect 125 1863 133 1864
rect 215 1863 223 1864
rect 125 1860 133 1861
rect 215 1860 223 1861
rect 2 1799 10 1800
rect 2 1796 10 1797
rect 24 1791 32 1792
rect 24 1788 32 1789
rect 88 1778 89 1786
rect 91 1778 92 1786
rect 107 1741 115 1742
rect 197 1741 205 1742
rect 107 1738 115 1739
rect 197 1738 205 1739
rect 129 1733 137 1734
rect 219 1733 227 1734
rect -165 1725 -164 1733
rect -162 1725 -161 1733
rect -126 1725 -125 1733
rect -123 1725 -122 1733
rect -86 1725 -85 1733
rect -83 1725 -82 1733
rect -47 1725 -46 1733
rect -44 1725 -43 1733
rect -6 1725 -5 1733
rect -3 1725 -2 1733
rect 129 1730 137 1731
rect 219 1730 227 1731
rect -177 1667 -176 1675
rect -174 1667 -173 1675
rect 103 1615 111 1616
rect 193 1615 201 1616
rect 103 1612 111 1613
rect 193 1612 201 1613
rect 125 1607 133 1608
rect 215 1607 223 1608
rect 125 1604 133 1605
rect 215 1604 223 1605
rect 2 1543 10 1544
rect 2 1540 10 1541
rect 24 1535 32 1536
rect 24 1532 32 1533
rect 88 1522 89 1530
rect 91 1522 92 1530
rect 1285 1516 1293 1517
rect 1375 1516 1383 1517
rect 1285 1513 1293 1514
rect 1375 1513 1383 1514
rect 1307 1508 1315 1509
rect 1397 1508 1405 1509
rect 324 1498 325 1506
rect 327 1498 328 1506
rect 1307 1505 1315 1506
rect 1397 1505 1405 1506
rect 107 1485 115 1486
rect 197 1485 205 1486
rect 107 1482 115 1483
rect 197 1482 205 1483
rect 359 1478 367 1479
rect 129 1477 137 1478
rect 219 1477 227 1478
rect -165 1469 -164 1477
rect -162 1469 -161 1477
rect -126 1469 -125 1477
rect -123 1469 -122 1477
rect -86 1469 -85 1477
rect -83 1469 -82 1477
rect -47 1469 -46 1477
rect -44 1469 -43 1477
rect -6 1469 -5 1477
rect -3 1469 -2 1477
rect 359 1475 367 1476
rect 129 1474 137 1475
rect 219 1474 227 1475
rect 381 1470 389 1471
rect 381 1467 389 1468
rect 1184 1444 1192 1445
rect 1184 1441 1192 1442
rect 445 1433 453 1434
rect 1206 1436 1214 1437
rect 325 1424 333 1425
rect 445 1430 453 1431
rect 467 1425 475 1426
rect 1206 1433 1214 1434
rect 325 1421 333 1422
rect -177 1411 -176 1419
rect -174 1411 -173 1419
rect 467 1422 475 1423
rect 1270 1423 1271 1431
rect 1273 1423 1274 1431
rect 359 1383 367 1384
rect 359 1380 367 1381
rect 1289 1386 1297 1387
rect 1379 1386 1387 1387
rect 1289 1383 1297 1384
rect 1379 1383 1387 1384
rect 1311 1378 1319 1379
rect 1401 1378 1409 1379
rect 381 1375 389 1376
rect 103 1359 111 1360
rect 193 1359 201 1360
rect 381 1372 389 1373
rect 1017 1370 1018 1378
rect 1020 1370 1021 1378
rect 1056 1370 1057 1378
rect 1059 1370 1060 1378
rect 1096 1370 1097 1378
rect 1099 1370 1100 1378
rect 1135 1370 1136 1378
rect 1138 1370 1139 1378
rect 1176 1370 1177 1378
rect 1179 1370 1180 1378
rect 1311 1375 1319 1376
rect 1401 1375 1409 1376
rect 103 1356 111 1357
rect 193 1356 201 1357
rect 784 1356 785 1364
rect 787 1356 788 1364
rect 125 1351 133 1352
rect 215 1351 223 1352
rect 125 1348 133 1349
rect 215 1348 223 1349
rect 819 1336 827 1337
rect 819 1333 827 1334
rect 841 1328 849 1329
rect 841 1325 849 1326
rect 1005 1312 1006 1320
rect 1008 1312 1009 1320
rect 2 1287 10 1288
rect 905 1291 913 1292
rect 2 1284 10 1285
rect 24 1279 32 1280
rect 24 1276 32 1277
rect 785 1282 793 1283
rect 905 1288 913 1289
rect 927 1283 935 1284
rect 88 1266 89 1274
rect 91 1266 92 1274
rect 314 1270 322 1271
rect 785 1279 793 1280
rect 927 1280 935 1281
rect 314 1267 322 1268
rect 336 1262 344 1263
rect 336 1259 344 1260
rect 401 1252 402 1260
rect 404 1252 405 1260
rect 1285 1260 1293 1261
rect 1375 1260 1383 1261
rect 1285 1257 1293 1258
rect 1375 1257 1383 1258
rect 1307 1252 1315 1253
rect 1397 1252 1405 1253
rect 819 1241 827 1242
rect 1307 1249 1315 1250
rect 1397 1249 1405 1250
rect 819 1238 827 1239
rect 107 1229 115 1230
rect 197 1229 205 1230
rect 841 1233 849 1234
rect 107 1226 115 1227
rect 197 1226 205 1227
rect 841 1230 849 1231
rect 129 1221 137 1222
rect 219 1221 227 1222
rect -165 1213 -164 1221
rect -162 1213 -161 1221
rect -126 1213 -125 1221
rect -123 1213 -122 1221
rect -86 1213 -85 1221
rect -83 1213 -82 1221
rect -47 1213 -46 1221
rect -44 1213 -43 1221
rect -6 1213 -5 1221
rect -3 1213 -2 1221
rect 129 1218 137 1219
rect 219 1218 227 1219
rect 1184 1188 1192 1189
rect 1184 1185 1192 1186
rect 1206 1180 1214 1181
rect 324 1163 325 1171
rect 327 1163 328 1171
rect 1206 1177 1214 1178
rect -177 1155 -176 1163
rect -174 1155 -173 1163
rect 1270 1167 1271 1175
rect 1273 1167 1274 1175
rect 359 1143 367 1144
rect 359 1140 367 1141
rect 381 1135 389 1136
rect 381 1132 389 1133
rect 784 1123 785 1131
rect 787 1123 788 1131
rect 1289 1130 1297 1131
rect 1379 1130 1387 1131
rect 1289 1127 1297 1128
rect 1379 1127 1387 1128
rect 1311 1122 1319 1123
rect 1401 1122 1409 1123
rect 1017 1114 1018 1122
rect 1020 1114 1021 1122
rect 1056 1114 1057 1122
rect 1059 1114 1060 1122
rect 1096 1114 1097 1122
rect 1099 1114 1100 1122
rect 1135 1114 1136 1122
rect 1138 1114 1139 1122
rect 1176 1114 1177 1122
rect 1179 1114 1180 1122
rect 1311 1119 1319 1120
rect 1401 1119 1409 1120
rect 103 1103 111 1104
rect 193 1103 201 1104
rect 103 1100 111 1101
rect 193 1100 201 1101
rect 445 1098 453 1099
rect 819 1103 827 1104
rect 819 1100 827 1101
rect 125 1095 133 1096
rect 215 1095 223 1096
rect 125 1092 133 1093
rect 215 1092 223 1093
rect 325 1089 333 1090
rect 445 1095 453 1096
rect 841 1095 849 1096
rect 467 1090 475 1091
rect 325 1086 333 1087
rect 467 1087 475 1088
rect 841 1092 849 1093
rect 905 1058 913 1059
rect 359 1048 367 1049
rect 785 1049 793 1050
rect 1005 1056 1006 1064
rect 1008 1056 1009 1064
rect 905 1055 913 1056
rect 927 1050 935 1051
rect 785 1046 793 1047
rect 359 1045 367 1046
rect 381 1040 389 1041
rect 927 1047 935 1048
rect 2 1031 10 1032
rect 2 1028 10 1029
rect 24 1023 32 1024
rect 24 1020 32 1021
rect 381 1037 389 1038
rect 88 1010 89 1018
rect 91 1010 92 1018
rect 729 1004 730 1012
rect 732 1004 733 1012
rect 819 1008 827 1009
rect 819 1005 827 1006
rect 1285 1004 1293 1005
rect 1375 1004 1383 1005
rect 841 1000 849 1001
rect 1285 1001 1293 1002
rect 1375 1001 1383 1002
rect 660 983 661 991
rect 663 983 664 991
rect 690 984 691 992
rect 693 984 694 992
rect 841 997 849 998
rect 1307 996 1315 997
rect 1397 996 1405 997
rect 1307 993 1315 994
rect 1397 993 1405 994
rect 107 973 115 974
rect 197 973 205 974
rect 107 970 115 971
rect 197 970 205 971
rect 129 965 137 966
rect 219 965 227 966
rect -165 957 -164 965
rect -162 957 -161 965
rect -126 957 -125 965
rect -123 957 -122 965
rect -86 957 -85 965
rect -83 957 -82 965
rect -47 957 -46 965
rect -44 957 -43 965
rect -6 957 -5 965
rect -3 957 -2 965
rect 129 962 137 963
rect 219 962 227 963
rect 652 953 653 961
rect 655 953 656 961
rect 314 935 322 936
rect 622 942 623 950
rect 625 942 626 950
rect 729 947 730 955
rect 732 947 733 955
rect 314 932 322 933
rect 336 927 344 928
rect 1184 932 1192 933
rect 336 924 344 925
rect 401 917 402 925
rect 404 917 405 925
rect 1184 929 1192 930
rect 1206 924 1214 925
rect 614 912 615 920
rect 617 912 618 920
rect 1206 921 1214 922
rect -177 899 -176 907
rect -174 899 -173 907
rect 584 901 585 909
rect 587 901 588 909
rect 1270 911 1271 919
rect 1273 911 1274 919
rect 729 890 730 898
rect 732 890 733 898
rect 784 890 785 898
rect 787 890 788 898
rect 576 871 577 879
rect 579 871 580 879
rect 819 870 827 871
rect 546 860 547 868
rect 549 860 550 868
rect 819 867 827 868
rect 1289 874 1297 875
rect 1379 874 1387 875
rect 1289 871 1297 872
rect 1379 871 1387 872
rect 1311 866 1319 867
rect 1401 866 1409 867
rect 841 862 849 863
rect 103 847 111 848
rect 193 847 201 848
rect 103 844 111 845
rect 193 844 201 845
rect 125 839 133 840
rect 215 839 223 840
rect 841 859 849 860
rect 1017 858 1018 866
rect 1020 858 1021 866
rect 1056 858 1057 866
rect 1059 858 1060 866
rect 1096 858 1097 866
rect 1099 858 1100 866
rect 1135 858 1136 866
rect 1138 858 1139 866
rect 1176 858 1177 866
rect 1179 858 1180 866
rect 1311 863 1319 864
rect 1401 863 1409 864
rect 125 836 133 837
rect 215 836 223 837
rect 324 828 325 836
rect 327 828 328 836
rect 538 831 539 839
rect 541 831 542 839
rect 729 833 730 841
rect 732 833 733 841
rect 905 825 913 826
rect 785 816 793 817
rect 905 822 913 823
rect 927 817 935 818
rect 359 808 367 809
rect 785 813 793 814
rect 359 805 367 806
rect 530 802 531 810
rect 533 802 534 810
rect 927 814 935 815
rect 381 800 389 801
rect 381 797 389 798
rect 1005 800 1006 808
rect 1008 800 1009 808
rect 2 775 10 776
rect 819 775 827 776
rect 2 772 10 773
rect 24 767 32 768
rect 24 764 32 765
rect 819 772 827 773
rect 445 763 453 764
rect 841 767 849 768
rect 88 754 89 762
rect 91 754 92 762
rect 325 754 333 755
rect 445 760 453 761
rect 841 764 849 765
rect 467 755 475 756
rect 325 751 333 752
rect 467 752 475 753
rect 1285 748 1293 749
rect 1375 748 1383 749
rect 1285 745 1293 746
rect 1375 745 1383 746
rect 1307 740 1315 741
rect 1397 740 1405 741
rect 1307 737 1315 738
rect 1397 737 1405 738
rect 107 717 115 718
rect 197 717 205 718
rect 107 714 115 715
rect 197 714 205 715
rect 359 713 367 714
rect 129 709 137 710
rect 219 709 227 710
rect 359 710 367 711
rect -165 701 -164 709
rect -162 701 -161 709
rect -126 701 -125 709
rect -123 701 -122 709
rect -86 701 -85 709
rect -83 701 -82 709
rect -47 701 -46 709
rect -44 701 -43 709
rect -6 701 -5 709
rect -3 701 -2 709
rect 129 706 137 707
rect 219 706 227 707
rect 381 705 389 706
rect 381 702 389 703
rect 1184 676 1192 677
rect 1184 673 1192 674
rect 1206 668 1214 669
rect 784 657 785 665
rect 787 657 788 665
rect 1206 665 1214 666
rect 1270 655 1271 663
rect 1273 655 1274 663
rect -177 643 -176 651
rect -174 643 -173 651
rect 819 637 827 638
rect 819 634 827 635
rect 841 629 849 630
rect 841 626 849 627
rect 1289 618 1297 619
rect 1379 618 1387 619
rect 1289 615 1297 616
rect 1379 615 1387 616
rect 1311 610 1319 611
rect 1401 610 1409 611
rect 314 600 322 601
rect 314 597 322 598
rect 103 591 111 592
rect 193 591 201 592
rect 336 592 344 593
rect 1017 602 1018 610
rect 1020 602 1021 610
rect 1056 602 1057 610
rect 1059 602 1060 610
rect 1096 602 1097 610
rect 1099 602 1100 610
rect 1135 602 1136 610
rect 1138 602 1139 610
rect 1176 602 1177 610
rect 1179 602 1180 610
rect 1311 607 1319 608
rect 1401 607 1409 608
rect 905 592 913 593
rect 103 588 111 589
rect 193 588 201 589
rect 125 583 133 584
rect 215 583 223 584
rect 336 589 344 590
rect 401 582 402 590
rect 404 582 405 590
rect 785 583 793 584
rect 905 589 913 590
rect 927 584 935 585
rect 125 580 133 581
rect 215 580 223 581
rect 785 580 793 581
rect 927 581 935 582
rect 819 542 827 543
rect 1005 544 1006 552
rect 1008 544 1009 552
rect 819 539 827 540
rect 841 534 849 535
rect 2 519 10 520
rect 841 531 849 532
rect 2 516 10 517
rect 24 511 32 512
rect 24 508 32 509
rect 88 498 89 506
rect 91 498 92 506
rect 324 493 325 501
rect 327 493 328 501
rect 1285 492 1293 493
rect 1375 492 1383 493
rect 1285 489 1293 490
rect 1375 489 1383 490
rect 784 481 785 489
rect 787 481 788 489
rect 1307 484 1315 485
rect 1397 484 1405 485
rect 359 473 367 474
rect 1307 481 1315 482
rect 1397 481 1405 482
rect 359 470 367 471
rect 107 461 115 462
rect 197 461 205 462
rect 381 465 389 466
rect 107 458 115 459
rect 197 458 205 459
rect 381 462 389 463
rect 129 453 137 454
rect 219 453 227 454
rect -165 445 -164 453
rect -162 445 -161 453
rect -126 445 -125 453
rect -123 445 -122 453
rect -86 445 -85 453
rect -83 445 -82 453
rect -47 445 -46 453
rect -44 445 -43 453
rect -6 445 -5 453
rect -3 445 -2 453
rect 129 450 137 451
rect 219 450 227 451
rect 445 428 453 429
rect 325 419 333 420
rect 445 425 453 426
rect 467 420 475 421
rect 1184 420 1192 421
rect 325 416 333 417
rect 467 417 475 418
rect 1184 417 1192 418
rect 1206 412 1214 413
rect 1206 409 1214 410
rect -177 387 -176 395
rect -174 387 -173 395
rect 1270 399 1271 407
rect 1273 399 1274 407
rect 359 378 367 379
rect 359 375 367 376
rect 381 370 389 371
rect 381 367 389 368
rect 1289 362 1297 363
rect 1379 362 1387 363
rect 1289 359 1297 360
rect 1379 359 1387 360
rect 1311 354 1319 355
rect 1401 354 1409 355
rect 1017 346 1018 354
rect 1020 346 1021 354
rect 1056 346 1057 354
rect 1059 346 1060 354
rect 1096 346 1097 354
rect 1099 346 1100 354
rect 1135 346 1136 354
rect 1138 346 1139 354
rect 1176 346 1177 354
rect 1179 346 1180 354
rect 1311 351 1319 352
rect 1401 351 1409 352
rect 103 335 111 336
rect 193 335 201 336
rect 103 332 111 333
rect 193 332 201 333
rect 125 327 133 328
rect 215 327 223 328
rect 125 324 133 325
rect 215 324 223 325
rect 1005 288 1006 296
rect 1008 288 1009 296
rect 2 263 10 264
rect 314 265 322 266
rect 314 262 322 263
rect 2 260 10 261
rect 24 255 32 256
rect 24 252 32 253
rect 336 257 344 258
rect 88 242 89 250
rect 91 242 92 250
rect 336 254 344 255
rect 401 247 402 255
rect 404 247 405 255
rect 107 205 115 206
rect 197 205 205 206
rect 107 202 115 203
rect 197 202 205 203
rect 129 197 137 198
rect 219 197 227 198
rect -165 189 -164 197
rect -162 189 -161 197
rect -126 189 -125 197
rect -123 189 -122 197
rect -86 189 -85 197
rect -83 189 -82 197
rect -47 189 -46 197
rect -44 189 -43 197
rect -6 189 -5 197
rect -3 189 -2 197
rect 129 194 137 195
rect 219 194 227 195
rect -177 131 -176 139
rect -174 131 -173 139
rect 103 79 111 80
rect 193 79 201 80
rect 103 76 111 77
rect 193 76 201 77
rect 125 71 133 72
rect 215 71 223 72
rect 125 68 133 69
rect 215 68 223 69
rect 2 7 10 8
rect 2 4 10 5
rect 24 -1 32 0
rect 24 -4 32 -3
rect 88 -14 89 -6
rect 91 -14 92 -6
rect 107 -51 115 -50
rect 197 -51 205 -50
rect 107 -54 115 -53
rect 197 -54 205 -53
rect 129 -59 137 -58
rect 219 -59 227 -58
rect -165 -67 -164 -59
rect -162 -67 -161 -59
rect -126 -67 -125 -59
rect -123 -67 -122 -59
rect -86 -67 -85 -59
rect -83 -67 -82 -59
rect -47 -67 -46 -59
rect -44 -67 -43 -59
rect -6 -67 -5 -59
rect -3 -67 -2 -59
rect 129 -62 137 -61
rect 219 -62 227 -61
rect -177 -125 -176 -117
rect -174 -125 -173 -117
<< pdiffusion >>
rect 149 1889 157 1890
rect 239 1889 247 1890
rect 149 1886 157 1887
rect 239 1886 247 1887
rect 149 1837 157 1838
rect 239 1837 247 1838
rect 149 1834 157 1835
rect 239 1834 247 1835
rect 48 1817 56 1818
rect 48 1814 56 1815
rect 88 1798 89 1806
rect 91 1798 92 1806
rect 48 1765 56 1766
rect 48 1762 56 1763
rect 153 1759 161 1760
rect 243 1759 251 1760
rect 153 1756 161 1757
rect -165 1745 -164 1753
rect -162 1745 -161 1753
rect -126 1745 -125 1753
rect -123 1745 -122 1753
rect -86 1745 -85 1753
rect -83 1745 -82 1753
rect -47 1745 -46 1753
rect -44 1745 -43 1753
rect -6 1745 -5 1753
rect -3 1745 -2 1753
rect 243 1756 251 1757
rect 153 1707 161 1708
rect 243 1707 251 1708
rect 153 1704 161 1705
rect 243 1704 251 1705
rect -177 1687 -176 1695
rect -174 1687 -173 1695
rect 149 1633 157 1634
rect 239 1633 247 1634
rect 149 1630 157 1631
rect 239 1630 247 1631
rect 149 1581 157 1582
rect 239 1581 247 1582
rect 149 1578 157 1579
rect 239 1578 247 1579
rect 48 1561 56 1562
rect 48 1558 56 1559
rect 88 1542 89 1550
rect 91 1542 92 1550
rect 1331 1534 1339 1535
rect 1421 1534 1429 1535
rect 1331 1531 1339 1532
rect 1421 1531 1429 1532
rect 324 1518 325 1526
rect 327 1518 328 1526
rect 48 1509 56 1510
rect 48 1506 56 1507
rect 153 1503 161 1504
rect 243 1503 251 1504
rect 153 1500 161 1501
rect -165 1489 -164 1497
rect -162 1489 -161 1497
rect -126 1489 -125 1497
rect -123 1489 -122 1497
rect -86 1489 -85 1497
rect -83 1489 -82 1497
rect -47 1489 -46 1497
rect -44 1489 -43 1497
rect -6 1489 -5 1497
rect -3 1489 -2 1497
rect 243 1500 251 1501
rect 405 1496 413 1497
rect 405 1493 413 1494
rect 1331 1482 1339 1483
rect 1421 1482 1429 1483
rect 1331 1479 1339 1480
rect 1421 1479 1429 1480
rect 1230 1462 1238 1463
rect 1230 1459 1238 1460
rect 153 1451 161 1452
rect 243 1451 251 1452
rect 491 1451 499 1452
rect 153 1448 161 1449
rect 243 1448 251 1449
rect 405 1444 413 1445
rect 491 1448 499 1449
rect -177 1431 -176 1439
rect -174 1431 -173 1439
rect 405 1441 413 1442
rect 1270 1443 1271 1451
rect 1273 1443 1274 1451
rect 345 1424 353 1425
rect 345 1421 353 1422
rect 1230 1410 1238 1411
rect 1230 1407 1238 1408
rect 405 1401 413 1402
rect 491 1399 499 1400
rect 405 1398 413 1399
rect 1335 1404 1343 1405
rect 1425 1404 1433 1405
rect 1335 1401 1343 1402
rect 491 1396 499 1397
rect 1017 1390 1018 1398
rect 1020 1390 1021 1398
rect 1056 1390 1057 1398
rect 1059 1390 1060 1398
rect 1096 1390 1097 1398
rect 1099 1390 1100 1398
rect 1135 1390 1136 1398
rect 1138 1390 1139 1398
rect 1176 1390 1177 1398
rect 1179 1390 1180 1398
rect 1425 1401 1433 1402
rect 149 1377 157 1378
rect 239 1377 247 1378
rect 784 1376 785 1384
rect 787 1376 788 1384
rect 149 1374 157 1375
rect 239 1374 247 1375
rect 865 1354 873 1355
rect 1335 1352 1343 1353
rect 1425 1352 1433 1353
rect 405 1349 413 1350
rect 865 1351 873 1352
rect 405 1346 413 1347
rect 1335 1349 1343 1350
rect 1425 1349 1433 1350
rect 149 1325 157 1326
rect 1005 1332 1006 1340
rect 1008 1332 1009 1340
rect 239 1325 247 1326
rect 149 1322 157 1323
rect 239 1322 247 1323
rect 951 1309 959 1310
rect 48 1305 56 1306
rect 48 1302 56 1303
rect 865 1302 873 1303
rect 951 1306 959 1307
rect 865 1299 873 1300
rect 88 1286 89 1294
rect 91 1286 92 1294
rect 360 1288 368 1289
rect 360 1285 368 1286
rect 805 1282 813 1283
rect 401 1272 402 1280
rect 404 1272 405 1280
rect 805 1279 813 1280
rect 1331 1278 1339 1279
rect 1421 1278 1429 1279
rect 1331 1275 1339 1276
rect 1421 1275 1429 1276
rect 48 1253 56 1254
rect 48 1250 56 1251
rect 153 1247 161 1248
rect 865 1259 873 1260
rect 951 1257 959 1258
rect 865 1256 873 1257
rect 243 1247 251 1248
rect 951 1254 959 1255
rect 153 1244 161 1245
rect -165 1233 -164 1241
rect -162 1233 -161 1241
rect -126 1233 -125 1241
rect -123 1233 -122 1241
rect -86 1233 -85 1241
rect -83 1233 -82 1241
rect -47 1233 -46 1241
rect -44 1233 -43 1241
rect -6 1233 -5 1241
rect -3 1233 -2 1241
rect 243 1244 251 1245
rect 360 1236 368 1237
rect 360 1233 368 1234
rect 1331 1226 1339 1227
rect 1421 1226 1429 1227
rect 1331 1223 1339 1224
rect 1421 1223 1429 1224
rect 865 1207 873 1208
rect 1230 1206 1238 1207
rect 865 1204 873 1205
rect 153 1195 161 1196
rect 1230 1203 1238 1204
rect 243 1195 251 1196
rect 153 1192 161 1193
rect 243 1192 251 1193
rect 324 1183 325 1191
rect 327 1183 328 1191
rect 1270 1187 1271 1195
rect 1273 1187 1274 1195
rect -177 1175 -176 1183
rect -174 1175 -173 1183
rect 405 1161 413 1162
rect 405 1158 413 1159
rect 1230 1154 1238 1155
rect 784 1143 785 1151
rect 787 1143 788 1151
rect 1230 1151 1238 1152
rect 149 1121 157 1122
rect 1335 1148 1343 1149
rect 1425 1148 1433 1149
rect 1335 1145 1343 1146
rect 1017 1134 1018 1142
rect 1020 1134 1021 1142
rect 1056 1134 1057 1142
rect 1059 1134 1060 1142
rect 1096 1134 1097 1142
rect 1099 1134 1100 1142
rect 1135 1134 1136 1142
rect 1138 1134 1139 1142
rect 1176 1134 1177 1142
rect 1179 1134 1180 1142
rect 1425 1145 1433 1146
rect 239 1121 247 1122
rect 149 1118 157 1119
rect 239 1118 247 1119
rect 865 1121 873 1122
rect 491 1116 499 1117
rect 865 1118 873 1119
rect 405 1109 413 1110
rect 491 1113 499 1114
rect 405 1106 413 1107
rect 1335 1096 1343 1097
rect 1425 1096 1433 1097
rect 345 1089 353 1090
rect 345 1086 353 1087
rect 1335 1093 1343 1094
rect 1425 1093 1433 1094
rect 951 1076 959 1077
rect 1005 1076 1006 1084
rect 1008 1076 1009 1084
rect 149 1069 157 1070
rect 239 1069 247 1070
rect 149 1066 157 1067
rect 239 1066 247 1067
rect 865 1069 873 1070
rect 951 1073 959 1074
rect 405 1066 413 1067
rect 491 1064 499 1065
rect 405 1063 413 1064
rect 865 1066 873 1067
rect 491 1061 499 1062
rect 48 1049 56 1050
rect 805 1049 813 1050
rect 48 1046 56 1047
rect 805 1046 813 1047
rect 88 1030 89 1038
rect 91 1030 92 1038
rect 546 1023 547 1031
rect 549 1023 550 1031
rect 584 1023 585 1031
rect 587 1023 588 1031
rect 622 1023 623 1031
rect 625 1023 626 1031
rect 660 1023 661 1031
rect 663 1023 664 1031
rect 729 1024 730 1032
rect 732 1024 733 1032
rect 865 1026 873 1027
rect 951 1024 959 1025
rect 405 1014 413 1015
rect 405 1011 413 1012
rect 865 1023 873 1024
rect 1331 1022 1339 1023
rect 1421 1022 1429 1023
rect 951 1021 959 1022
rect 1331 1019 1339 1020
rect 1421 1019 1429 1020
rect 48 997 56 998
rect 48 994 56 995
rect 153 991 161 992
rect 243 991 251 992
rect 153 988 161 989
rect -165 977 -164 985
rect -162 977 -161 985
rect -126 977 -125 985
rect -123 977 -122 985
rect -86 977 -85 985
rect -83 977 -82 985
rect -47 977 -46 985
rect -44 977 -43 985
rect -6 977 -5 985
rect -3 977 -2 985
rect 243 988 251 989
rect 729 967 730 975
rect 732 967 733 975
rect 865 974 873 975
rect 865 971 873 972
rect 360 953 368 954
rect 1331 970 1339 971
rect 1421 970 1429 971
rect 1331 967 1339 968
rect 1421 967 1429 968
rect 360 950 368 951
rect 153 939 161 940
rect 243 939 251 940
rect 153 936 161 937
rect 243 936 251 937
rect 401 937 402 945
rect 404 937 405 945
rect 1230 950 1238 951
rect 1230 947 1238 948
rect -177 919 -176 927
rect -174 919 -173 927
rect 1270 931 1271 939
rect 1273 931 1274 939
rect 729 910 730 918
rect 732 910 733 918
rect 784 910 785 918
rect 787 910 788 918
rect 360 901 368 902
rect 360 898 368 899
rect 1230 898 1238 899
rect 1230 895 1238 896
rect 865 888 873 889
rect 1335 892 1343 893
rect 1425 892 1433 893
rect 1335 889 1343 890
rect 865 885 873 886
rect 149 865 157 866
rect 1017 878 1018 886
rect 1020 878 1021 886
rect 1056 878 1057 886
rect 1059 878 1060 886
rect 1096 878 1097 886
rect 1099 878 1100 886
rect 1135 878 1136 886
rect 1138 878 1139 886
rect 1176 878 1177 886
rect 1179 878 1180 886
rect 1425 889 1433 890
rect 239 865 247 866
rect 149 862 157 863
rect 239 862 247 863
rect 324 848 325 856
rect 327 848 328 856
rect 729 853 730 861
rect 732 853 733 861
rect 951 843 959 844
rect 865 836 873 837
rect 951 840 959 841
rect 1335 840 1343 841
rect 1425 840 1433 841
rect 865 833 873 834
rect 405 826 413 827
rect 1335 837 1343 838
rect 1425 837 1433 838
rect 405 823 413 824
rect 149 813 157 814
rect 1005 820 1006 828
rect 1008 820 1009 828
rect 805 816 813 817
rect 239 813 247 814
rect 149 810 157 811
rect 239 810 247 811
rect 805 813 813 814
rect 48 793 56 794
rect 48 790 56 791
rect 865 793 873 794
rect 951 791 959 792
rect 865 790 873 791
rect 88 774 89 782
rect 91 774 92 782
rect 951 788 959 789
rect 491 781 499 782
rect 405 774 413 775
rect 491 778 499 779
rect 405 771 413 772
rect 1331 766 1339 767
rect 1421 766 1429 767
rect 1331 763 1339 764
rect 1421 763 1429 764
rect 345 754 353 755
rect 345 751 353 752
rect 48 741 56 742
rect 48 738 56 739
rect 865 741 873 742
rect 153 735 161 736
rect 243 735 251 736
rect 153 732 161 733
rect -165 721 -164 729
rect -162 721 -161 729
rect -126 721 -125 729
rect -123 721 -122 729
rect -86 721 -85 729
rect -83 721 -82 729
rect -47 721 -46 729
rect -44 721 -43 729
rect -6 721 -5 729
rect -3 721 -2 729
rect 243 732 251 733
rect 865 738 873 739
rect 405 731 413 732
rect 491 729 499 730
rect 405 728 413 729
rect 491 726 499 727
rect 1331 714 1339 715
rect 1421 714 1429 715
rect 1331 711 1339 712
rect 1421 711 1429 712
rect 1230 694 1238 695
rect 1230 691 1238 692
rect 153 683 161 684
rect 243 683 251 684
rect 153 680 161 681
rect 243 680 251 681
rect 405 679 413 680
rect 784 677 785 685
rect 787 677 788 685
rect 405 676 413 677
rect -177 663 -176 671
rect -174 663 -173 671
rect 1270 675 1271 683
rect 1273 675 1274 683
rect 865 655 873 656
rect 865 652 873 653
rect 1230 642 1238 643
rect 1230 639 1238 640
rect 1335 636 1343 637
rect 1425 636 1433 637
rect 1335 633 1343 634
rect 360 618 368 619
rect 1017 622 1018 630
rect 1020 622 1021 630
rect 1056 622 1057 630
rect 1059 622 1060 630
rect 1096 622 1097 630
rect 1099 622 1100 630
rect 1135 622 1136 630
rect 1138 622 1139 630
rect 1176 622 1177 630
rect 1179 622 1180 630
rect 1425 633 1433 634
rect 360 615 368 616
rect 149 609 157 610
rect 951 610 959 611
rect 239 609 247 610
rect 149 606 157 607
rect 239 606 247 607
rect 401 602 402 610
rect 404 602 405 610
rect 865 603 873 604
rect 951 607 959 608
rect 865 600 873 601
rect 1335 584 1343 585
rect 1425 584 1433 585
rect 805 583 813 584
rect 805 580 813 581
rect 1335 581 1343 582
rect 1425 581 1433 582
rect 360 566 368 567
rect 149 557 157 558
rect 360 563 368 564
rect 239 557 247 558
rect 1005 564 1006 572
rect 1008 564 1009 572
rect 865 560 873 561
rect 951 558 959 559
rect 865 557 873 558
rect 149 554 157 555
rect 239 554 247 555
rect 951 555 959 556
rect 48 537 56 538
rect 48 534 56 535
rect 88 518 89 526
rect 91 518 92 526
rect 324 513 325 521
rect 327 513 328 521
rect 1331 510 1339 511
rect 1421 510 1429 511
rect 784 501 785 509
rect 787 501 788 509
rect 865 508 873 509
rect 1331 507 1339 508
rect 865 505 873 506
rect 405 491 413 492
rect 1421 507 1429 508
rect 405 488 413 489
rect 48 485 56 486
rect 48 482 56 483
rect 153 479 161 480
rect 243 479 251 480
rect 153 476 161 477
rect -165 465 -164 473
rect -162 465 -161 473
rect -126 465 -125 473
rect -123 465 -122 473
rect -86 465 -85 473
rect -83 465 -82 473
rect -47 465 -46 473
rect -44 465 -43 473
rect -6 465 -5 473
rect -3 465 -2 473
rect 243 476 251 477
rect 1331 458 1339 459
rect 1421 458 1429 459
rect 1331 455 1339 456
rect 1421 455 1429 456
rect 491 446 499 447
rect 405 439 413 440
rect 491 443 499 444
rect 1230 438 1238 439
rect 405 436 413 437
rect 153 427 161 428
rect 243 427 251 428
rect 1230 435 1238 436
rect 153 424 161 425
rect 243 424 251 425
rect 345 419 353 420
rect 1270 419 1271 427
rect 1273 419 1274 427
rect -177 407 -176 415
rect -174 407 -173 415
rect 345 416 353 417
rect 405 396 413 397
rect 491 394 499 395
rect 405 393 413 394
rect 491 391 499 392
rect 1230 386 1238 387
rect 1230 383 1238 384
rect 1335 380 1343 381
rect 1425 380 1433 381
rect 1335 377 1343 378
rect 1017 366 1018 374
rect 1020 366 1021 374
rect 1056 366 1057 374
rect 1059 366 1060 374
rect 1096 366 1097 374
rect 1099 366 1100 374
rect 1135 366 1136 374
rect 1138 366 1139 374
rect 1176 366 1177 374
rect 1179 366 1180 374
rect 1425 377 1433 378
rect 149 353 157 354
rect 239 353 247 354
rect 149 350 157 351
rect 239 350 247 351
rect 405 344 413 345
rect 405 341 413 342
rect 1335 328 1343 329
rect 1425 328 1433 329
rect 1335 325 1343 326
rect 1425 325 1433 326
rect 1005 308 1006 316
rect 1008 308 1009 316
rect 149 301 157 302
rect 239 301 247 302
rect 149 298 157 299
rect 239 298 247 299
rect 360 283 368 284
rect 48 281 56 282
rect 360 280 368 281
rect 48 278 56 279
rect 88 262 89 270
rect 91 262 92 270
rect 401 267 402 275
rect 404 267 405 275
rect 360 231 368 232
rect 48 229 56 230
rect 48 226 56 227
rect 153 223 161 224
rect 360 228 368 229
rect 243 223 251 224
rect 153 220 161 221
rect -165 209 -164 217
rect -162 209 -161 217
rect -126 209 -125 217
rect -123 209 -122 217
rect -86 209 -85 217
rect -83 209 -82 217
rect -47 209 -46 217
rect -44 209 -43 217
rect -6 209 -5 217
rect -3 209 -2 217
rect 243 220 251 221
rect 153 171 161 172
rect 243 171 251 172
rect 153 168 161 169
rect 243 168 251 169
rect -177 151 -176 159
rect -174 151 -173 159
rect 149 97 157 98
rect 239 97 247 98
rect 149 94 157 95
rect 239 94 247 95
rect 149 45 157 46
rect 239 45 247 46
rect 149 42 157 43
rect 239 42 247 43
rect 48 25 56 26
rect 48 22 56 23
rect 88 6 89 14
rect 91 6 92 14
rect 48 -27 56 -26
rect 48 -30 56 -29
rect 153 -33 161 -32
rect 243 -33 251 -32
rect 153 -36 161 -35
rect -165 -47 -164 -39
rect -162 -47 -161 -39
rect -126 -47 -125 -39
rect -123 -47 -122 -39
rect -86 -47 -85 -39
rect -83 -47 -82 -39
rect -47 -47 -46 -39
rect -44 -47 -43 -39
rect -6 -47 -5 -39
rect -3 -47 -2 -39
rect 243 -36 251 -35
rect 153 -85 161 -84
rect 243 -85 251 -84
rect 153 -88 161 -87
rect 243 -88 251 -87
rect -177 -105 -176 -97
rect -174 -105 -173 -97
<< ndcontact >>
rect 103 1872 111 1876
rect 193 1872 201 1876
rect 103 1864 111 1868
rect 125 1864 133 1868
rect 193 1864 201 1868
rect 215 1864 223 1868
rect 125 1856 133 1860
rect 215 1856 223 1860
rect 2 1800 10 1804
rect 2 1792 10 1796
rect 24 1792 32 1796
rect 24 1784 32 1788
rect 84 1778 88 1786
rect 92 1778 96 1786
rect 107 1742 115 1746
rect 197 1742 205 1746
rect 107 1734 115 1738
rect 129 1734 137 1738
rect 197 1734 205 1738
rect 219 1734 227 1738
rect -169 1725 -165 1733
rect -161 1725 -157 1733
rect -130 1725 -126 1733
rect -122 1725 -118 1733
rect -90 1725 -86 1733
rect -82 1725 -78 1733
rect -51 1725 -47 1733
rect -43 1725 -39 1733
rect -10 1725 -6 1733
rect -2 1725 2 1733
rect 129 1726 137 1730
rect 219 1726 227 1730
rect -181 1667 -177 1675
rect -173 1667 -169 1675
rect 103 1616 111 1620
rect 193 1616 201 1620
rect 103 1608 111 1612
rect 125 1608 133 1612
rect 193 1608 201 1612
rect 215 1608 223 1612
rect 125 1600 133 1604
rect 215 1600 223 1604
rect 2 1544 10 1548
rect 2 1536 10 1540
rect 24 1536 32 1540
rect 24 1528 32 1532
rect 84 1522 88 1530
rect 92 1522 96 1530
rect 1285 1517 1293 1521
rect 1375 1517 1383 1521
rect 1285 1509 1293 1513
rect 1307 1509 1315 1513
rect 1375 1509 1383 1513
rect 1397 1509 1405 1513
rect 320 1498 324 1506
rect 328 1498 332 1506
rect 1307 1501 1315 1505
rect 1397 1501 1405 1505
rect 107 1486 115 1490
rect 197 1486 205 1490
rect 107 1478 115 1482
rect 129 1478 137 1482
rect 197 1478 205 1482
rect 219 1478 227 1482
rect 359 1479 367 1483
rect -169 1469 -165 1477
rect -161 1469 -157 1477
rect -130 1469 -126 1477
rect -122 1469 -118 1477
rect -90 1469 -86 1477
rect -82 1469 -78 1477
rect -51 1469 -47 1477
rect -43 1469 -39 1477
rect -10 1469 -6 1477
rect -2 1469 2 1477
rect 129 1470 137 1474
rect 219 1470 227 1474
rect 359 1471 367 1475
rect 381 1471 389 1475
rect 381 1463 389 1467
rect 1184 1445 1192 1449
rect 445 1434 453 1438
rect 1184 1437 1192 1441
rect 1206 1437 1214 1441
rect 325 1425 333 1429
rect 445 1426 453 1430
rect 467 1426 475 1430
rect 1206 1429 1214 1433
rect -181 1411 -177 1419
rect -173 1411 -169 1419
rect 325 1417 333 1421
rect 467 1418 475 1422
rect 1266 1423 1270 1431
rect 1274 1423 1278 1431
rect 359 1384 367 1388
rect 359 1376 367 1380
rect 381 1376 389 1380
rect 1289 1387 1297 1391
rect 1379 1387 1387 1391
rect 1289 1379 1297 1383
rect 1311 1379 1319 1383
rect 1379 1379 1387 1383
rect 1401 1379 1409 1383
rect 103 1360 111 1364
rect 193 1360 201 1364
rect 381 1368 389 1372
rect 1013 1370 1017 1378
rect 1021 1370 1025 1378
rect 1052 1370 1056 1378
rect 1060 1370 1064 1378
rect 1092 1370 1096 1378
rect 1100 1370 1104 1378
rect 1131 1370 1135 1378
rect 1139 1370 1143 1378
rect 1172 1370 1176 1378
rect 1180 1370 1184 1378
rect 1311 1371 1319 1375
rect 1401 1371 1409 1375
rect 780 1356 784 1364
rect 788 1356 792 1364
rect 103 1352 111 1356
rect 125 1352 133 1356
rect 193 1352 201 1356
rect 215 1352 223 1356
rect 125 1344 133 1348
rect 215 1344 223 1348
rect 819 1337 827 1341
rect 819 1329 827 1333
rect 841 1329 849 1333
rect 841 1321 849 1325
rect 1001 1312 1005 1320
rect 1009 1312 1013 1320
rect 2 1288 10 1292
rect 905 1292 913 1296
rect 2 1280 10 1284
rect 24 1280 32 1284
rect 24 1272 32 1276
rect 785 1283 793 1287
rect 905 1284 913 1288
rect 927 1284 935 1288
rect 84 1266 88 1274
rect 92 1266 96 1274
rect 314 1271 322 1275
rect 785 1275 793 1279
rect 927 1276 935 1280
rect 314 1263 322 1267
rect 336 1263 344 1267
rect 336 1255 344 1259
rect 397 1252 401 1260
rect 405 1252 409 1260
rect 1285 1261 1293 1265
rect 1375 1261 1383 1265
rect 1285 1253 1293 1257
rect 1307 1253 1315 1257
rect 1375 1253 1383 1257
rect 1397 1253 1405 1257
rect 819 1242 827 1246
rect 1307 1245 1315 1249
rect 1397 1245 1405 1249
rect 107 1230 115 1234
rect 197 1230 205 1234
rect 819 1234 827 1238
rect 841 1234 849 1238
rect 107 1222 115 1226
rect 129 1222 137 1226
rect 197 1222 205 1226
rect 219 1222 227 1226
rect 841 1226 849 1230
rect -169 1213 -165 1221
rect -161 1213 -157 1221
rect -130 1213 -126 1221
rect -122 1213 -118 1221
rect -90 1213 -86 1221
rect -82 1213 -78 1221
rect -51 1213 -47 1221
rect -43 1213 -39 1221
rect -10 1213 -6 1221
rect -2 1213 2 1221
rect 129 1214 137 1218
rect 219 1214 227 1218
rect 1184 1189 1192 1193
rect 1184 1181 1192 1185
rect 1206 1181 1214 1185
rect 320 1163 324 1171
rect 328 1163 332 1171
rect 1206 1173 1214 1177
rect -181 1155 -177 1163
rect -173 1155 -169 1163
rect 1266 1167 1270 1175
rect 1274 1167 1278 1175
rect 359 1144 367 1148
rect 359 1136 367 1140
rect 381 1136 389 1140
rect 381 1128 389 1132
rect 780 1123 784 1131
rect 788 1123 792 1131
rect 1289 1131 1297 1135
rect 1379 1131 1387 1135
rect 1289 1123 1297 1127
rect 1311 1123 1319 1127
rect 1379 1123 1387 1127
rect 1401 1123 1409 1127
rect 1013 1114 1017 1122
rect 1021 1114 1025 1122
rect 1052 1114 1056 1122
rect 1060 1114 1064 1122
rect 1092 1114 1096 1122
rect 1100 1114 1104 1122
rect 1131 1114 1135 1122
rect 1139 1114 1143 1122
rect 1172 1114 1176 1122
rect 1180 1114 1184 1122
rect 1311 1115 1319 1119
rect 1401 1115 1409 1119
rect 103 1104 111 1108
rect 193 1104 201 1108
rect 103 1096 111 1100
rect 125 1096 133 1100
rect 193 1096 201 1100
rect 215 1096 223 1100
rect 819 1104 827 1108
rect 445 1099 453 1103
rect 125 1088 133 1092
rect 215 1088 223 1092
rect 325 1090 333 1094
rect 819 1096 827 1100
rect 841 1096 849 1100
rect 445 1091 453 1095
rect 467 1091 475 1095
rect 325 1082 333 1086
rect 467 1083 475 1087
rect 841 1088 849 1092
rect 905 1059 913 1063
rect 359 1049 367 1053
rect 785 1050 793 1054
rect 1001 1056 1005 1064
rect 1009 1056 1013 1064
rect 905 1051 913 1055
rect 927 1051 935 1055
rect 359 1041 367 1045
rect 381 1041 389 1045
rect 785 1042 793 1046
rect 927 1043 935 1047
rect 2 1032 10 1036
rect 2 1024 10 1028
rect 24 1024 32 1028
rect 24 1016 32 1020
rect 381 1033 389 1037
rect 84 1010 88 1018
rect 92 1010 96 1018
rect 725 1004 729 1012
rect 733 1004 737 1012
rect 819 1009 827 1013
rect 1285 1005 1293 1009
rect 819 1001 827 1005
rect 841 1001 849 1005
rect 1375 1005 1383 1009
rect 656 983 660 991
rect 664 983 668 991
rect 686 984 690 992
rect 694 984 698 992
rect 1285 997 1293 1001
rect 1307 997 1315 1001
rect 1375 997 1383 1001
rect 1397 997 1405 1001
rect 841 993 849 997
rect 1307 989 1315 993
rect 1397 989 1405 993
rect 107 974 115 978
rect 197 974 205 978
rect 107 966 115 970
rect 129 966 137 970
rect 197 966 205 970
rect 219 966 227 970
rect -169 957 -165 965
rect -161 957 -157 965
rect -130 957 -126 965
rect -122 957 -118 965
rect -90 957 -86 965
rect -82 957 -78 965
rect -51 957 -47 965
rect -43 957 -39 965
rect -10 957 -6 965
rect -2 957 2 965
rect 129 958 137 962
rect 219 958 227 962
rect 648 953 652 961
rect 656 953 660 961
rect 314 936 322 940
rect 618 942 622 950
rect 626 942 630 950
rect 725 947 729 955
rect 733 947 737 955
rect 314 928 322 932
rect 336 928 344 932
rect 1184 933 1192 937
rect 336 920 344 924
rect 397 917 401 925
rect 405 917 409 925
rect 1184 925 1192 929
rect 1206 925 1214 929
rect 610 912 614 920
rect 618 912 622 920
rect 1206 917 1214 921
rect -181 899 -177 907
rect -173 899 -169 907
rect 580 901 584 909
rect 588 901 592 909
rect 1266 911 1270 919
rect 1274 911 1278 919
rect 725 890 729 898
rect 733 890 737 898
rect 780 890 784 898
rect 788 890 792 898
rect 572 871 576 879
rect 580 871 584 879
rect 819 871 827 875
rect 542 860 546 868
rect 550 860 554 868
rect 819 863 827 867
rect 841 863 849 867
rect 1289 875 1297 879
rect 1379 875 1387 879
rect 1289 867 1297 871
rect 1311 867 1319 871
rect 1379 867 1387 871
rect 1401 867 1409 871
rect 103 848 111 852
rect 193 848 201 852
rect 103 840 111 844
rect 125 840 133 844
rect 193 840 201 844
rect 215 840 223 844
rect 841 855 849 859
rect 1013 858 1017 866
rect 1021 858 1025 866
rect 1052 858 1056 866
rect 1060 858 1064 866
rect 1092 858 1096 866
rect 1100 858 1104 866
rect 1131 858 1135 866
rect 1139 858 1143 866
rect 1172 858 1176 866
rect 1180 858 1184 866
rect 1311 859 1319 863
rect 1401 859 1409 863
rect 125 832 133 836
rect 215 832 223 836
rect 320 828 324 836
rect 328 828 332 836
rect 534 831 538 839
rect 542 831 546 839
rect 725 833 729 841
rect 733 833 737 841
rect 905 826 913 830
rect 785 817 793 821
rect 905 818 913 822
rect 927 818 935 822
rect 359 809 367 813
rect 359 801 367 805
rect 381 801 389 805
rect 526 802 530 810
rect 534 802 538 810
rect 785 809 793 813
rect 927 810 935 814
rect 1001 800 1005 808
rect 1009 800 1013 808
rect 381 793 389 797
rect 2 776 10 780
rect 819 776 827 780
rect 2 768 10 772
rect 24 768 32 772
rect 24 760 32 764
rect 445 764 453 768
rect 819 768 827 772
rect 841 768 849 772
rect 84 754 88 762
rect 92 754 96 762
rect 325 755 333 759
rect 445 756 453 760
rect 467 756 475 760
rect 841 760 849 764
rect 325 747 333 751
rect 467 748 475 752
rect 1285 749 1293 753
rect 1375 749 1383 753
rect 1285 741 1293 745
rect 1307 741 1315 745
rect 1375 741 1383 745
rect 1397 741 1405 745
rect 1307 733 1315 737
rect 1397 733 1405 737
rect 107 718 115 722
rect 197 718 205 722
rect 359 714 367 718
rect 107 710 115 714
rect 129 710 137 714
rect 197 710 205 714
rect 219 710 227 714
rect -169 701 -165 709
rect -161 701 -157 709
rect -130 701 -126 709
rect -122 701 -118 709
rect -90 701 -86 709
rect -82 701 -78 709
rect -51 701 -47 709
rect -43 701 -39 709
rect -10 701 -6 709
rect -2 701 2 709
rect 129 702 137 706
rect 359 706 367 710
rect 381 706 389 710
rect 219 702 227 706
rect 381 698 389 702
rect 1184 677 1192 681
rect 1184 669 1192 673
rect 1206 669 1214 673
rect 780 657 784 665
rect 788 657 792 665
rect 1206 661 1214 665
rect 1266 655 1270 663
rect 1274 655 1278 663
rect -181 643 -177 651
rect -173 643 -169 651
rect 819 638 827 642
rect 819 630 827 634
rect 841 630 849 634
rect 841 622 849 626
rect 1289 619 1297 623
rect 1379 619 1387 623
rect 1289 611 1297 615
rect 1311 611 1319 615
rect 1379 611 1387 615
rect 1401 611 1409 615
rect 314 601 322 605
rect 103 592 111 596
rect 193 592 201 596
rect 314 593 322 597
rect 336 593 344 597
rect 1013 602 1017 610
rect 1021 602 1025 610
rect 1052 602 1056 610
rect 1060 602 1064 610
rect 1092 602 1096 610
rect 1100 602 1104 610
rect 1131 602 1135 610
rect 1139 602 1143 610
rect 1172 602 1176 610
rect 1180 602 1184 610
rect 1311 603 1319 607
rect 1401 603 1409 607
rect 905 593 913 597
rect 103 584 111 588
rect 125 584 133 588
rect 193 584 201 588
rect 215 584 223 588
rect 336 585 344 589
rect 397 582 401 590
rect 405 582 409 590
rect 785 584 793 588
rect 905 585 913 589
rect 927 585 935 589
rect 125 576 133 580
rect 215 576 223 580
rect 785 576 793 580
rect 927 577 935 581
rect 819 543 827 547
rect 1001 544 1005 552
rect 1009 544 1013 552
rect 819 535 827 539
rect 841 535 849 539
rect 2 520 10 524
rect 841 527 849 531
rect 2 512 10 516
rect 24 512 32 516
rect 24 504 32 508
rect 84 498 88 506
rect 92 498 96 506
rect 320 493 324 501
rect 328 493 332 501
rect 1285 493 1293 497
rect 1375 493 1383 497
rect 780 481 784 489
rect 788 481 792 489
rect 1285 485 1293 489
rect 1307 485 1315 489
rect 1375 485 1383 489
rect 1397 485 1405 489
rect 359 474 367 478
rect 1307 477 1315 481
rect 1397 477 1405 481
rect 107 462 115 466
rect 197 462 205 466
rect 359 466 367 470
rect 381 466 389 470
rect 107 454 115 458
rect 129 454 137 458
rect 197 454 205 458
rect 219 454 227 458
rect 381 458 389 462
rect -169 445 -165 453
rect -161 445 -157 453
rect -130 445 -126 453
rect -122 445 -118 453
rect -90 445 -86 453
rect -82 445 -78 453
rect -51 445 -47 453
rect -43 445 -39 453
rect -10 445 -6 453
rect -2 445 2 453
rect 129 446 137 450
rect 219 446 227 450
rect 445 429 453 433
rect 325 420 333 424
rect 445 421 453 425
rect 467 421 475 425
rect 1184 421 1192 425
rect 325 412 333 416
rect 467 413 475 417
rect 1184 413 1192 417
rect 1206 413 1214 417
rect 1206 405 1214 409
rect -181 387 -177 395
rect -173 387 -169 395
rect 1266 399 1270 407
rect 1274 399 1278 407
rect 359 379 367 383
rect 359 371 367 375
rect 381 371 389 375
rect 381 363 389 367
rect 1289 363 1297 367
rect 1379 363 1387 367
rect 1289 355 1297 359
rect 1311 355 1319 359
rect 1379 355 1387 359
rect 1401 355 1409 359
rect 1013 346 1017 354
rect 1021 346 1025 354
rect 1052 346 1056 354
rect 1060 346 1064 354
rect 1092 346 1096 354
rect 1100 346 1104 354
rect 1131 346 1135 354
rect 1139 346 1143 354
rect 1172 346 1176 354
rect 1180 346 1184 354
rect 1311 347 1319 351
rect 1401 347 1409 351
rect 103 336 111 340
rect 193 336 201 340
rect 103 328 111 332
rect 125 328 133 332
rect 193 328 201 332
rect 215 328 223 332
rect 125 320 133 324
rect 215 320 223 324
rect 1001 288 1005 296
rect 1009 288 1013 296
rect 2 264 10 268
rect 314 266 322 270
rect 2 256 10 260
rect 24 256 32 260
rect 24 248 32 252
rect 314 258 322 262
rect 336 258 344 262
rect 84 242 88 250
rect 92 242 96 250
rect 336 250 344 254
rect 397 247 401 255
rect 405 247 409 255
rect 107 206 115 210
rect 197 206 205 210
rect 107 198 115 202
rect 129 198 137 202
rect 197 198 205 202
rect 219 198 227 202
rect -169 189 -165 197
rect -161 189 -157 197
rect -130 189 -126 197
rect -122 189 -118 197
rect -90 189 -86 197
rect -82 189 -78 197
rect -51 189 -47 197
rect -43 189 -39 197
rect -10 189 -6 197
rect -2 189 2 197
rect 129 190 137 194
rect 219 190 227 194
rect -181 131 -177 139
rect -173 131 -169 139
rect 103 80 111 84
rect 193 80 201 84
rect 103 72 111 76
rect 125 72 133 76
rect 193 72 201 76
rect 215 72 223 76
rect 125 64 133 68
rect 215 64 223 68
rect 2 8 10 12
rect 2 0 10 4
rect 24 0 32 4
rect 24 -8 32 -4
rect 84 -14 88 -6
rect 92 -14 96 -6
rect 107 -50 115 -46
rect 197 -50 205 -46
rect 107 -58 115 -54
rect 129 -58 137 -54
rect 197 -58 205 -54
rect 219 -58 227 -54
rect -169 -67 -165 -59
rect -161 -67 -157 -59
rect -130 -67 -126 -59
rect -122 -67 -118 -59
rect -90 -67 -86 -59
rect -82 -67 -78 -59
rect -51 -67 -47 -59
rect -43 -67 -39 -59
rect -10 -67 -6 -59
rect -2 -67 2 -59
rect 129 -66 137 -62
rect 219 -66 227 -62
rect -181 -125 -177 -117
rect -173 -125 -169 -117
<< pdcontact >>
rect 149 1890 157 1894
rect 239 1890 247 1894
rect 149 1882 157 1886
rect 239 1882 247 1886
rect 149 1838 157 1842
rect 239 1838 247 1842
rect 149 1830 157 1834
rect 239 1830 247 1834
rect 48 1818 56 1822
rect 48 1810 56 1814
rect 84 1798 88 1806
rect 92 1798 96 1806
rect 48 1766 56 1770
rect 48 1758 56 1762
rect 153 1760 161 1764
rect 243 1760 251 1764
rect -169 1745 -165 1753
rect -161 1745 -157 1753
rect -130 1745 -126 1753
rect -122 1745 -118 1753
rect -90 1745 -86 1753
rect -82 1745 -78 1753
rect -51 1745 -47 1753
rect -43 1745 -39 1753
rect -10 1745 -6 1753
rect -2 1745 2 1753
rect 153 1752 161 1756
rect 243 1752 251 1756
rect 153 1708 161 1712
rect 243 1708 251 1712
rect 153 1700 161 1704
rect 243 1700 251 1704
rect -181 1687 -177 1695
rect -173 1687 -169 1695
rect 149 1634 157 1638
rect 239 1634 247 1638
rect 149 1626 157 1630
rect 239 1626 247 1630
rect 149 1582 157 1586
rect 239 1582 247 1586
rect 149 1574 157 1578
rect 239 1574 247 1578
rect 48 1562 56 1566
rect 48 1554 56 1558
rect 84 1542 88 1550
rect 92 1542 96 1550
rect 1331 1535 1339 1539
rect 1421 1535 1429 1539
rect 1331 1527 1339 1531
rect 1421 1527 1429 1531
rect 320 1518 324 1526
rect 328 1518 332 1526
rect 48 1510 56 1514
rect 48 1502 56 1506
rect 153 1504 161 1508
rect 243 1504 251 1508
rect -169 1489 -165 1497
rect -161 1489 -157 1497
rect -130 1489 -126 1497
rect -122 1489 -118 1497
rect -90 1489 -86 1497
rect -82 1489 -78 1497
rect -51 1489 -47 1497
rect -43 1489 -39 1497
rect -10 1489 -6 1497
rect -2 1489 2 1497
rect 153 1496 161 1500
rect 243 1496 251 1500
rect 405 1497 413 1501
rect 405 1489 413 1493
rect 1331 1483 1339 1487
rect 1421 1483 1429 1487
rect 1331 1475 1339 1479
rect 1421 1475 1429 1479
rect 1230 1463 1238 1467
rect 153 1452 161 1456
rect 243 1452 251 1456
rect 491 1452 499 1456
rect 1230 1455 1238 1459
rect 153 1444 161 1448
rect 243 1444 251 1448
rect 405 1445 413 1449
rect 491 1444 499 1448
rect -181 1431 -177 1439
rect -173 1431 -169 1439
rect 405 1437 413 1441
rect 1266 1443 1270 1451
rect 1274 1443 1278 1451
rect 345 1425 353 1429
rect 345 1417 353 1421
rect 1230 1411 1238 1415
rect 405 1402 413 1406
rect 491 1400 499 1404
rect 405 1394 413 1398
rect 1230 1403 1238 1407
rect 1335 1405 1343 1409
rect 1425 1405 1433 1409
rect 491 1392 499 1396
rect 1013 1390 1017 1398
rect 1021 1390 1025 1398
rect 1052 1390 1056 1398
rect 1060 1390 1064 1398
rect 1092 1390 1096 1398
rect 1100 1390 1104 1398
rect 1131 1390 1135 1398
rect 1139 1390 1143 1398
rect 1172 1390 1176 1398
rect 1180 1390 1184 1398
rect 1335 1397 1343 1401
rect 1425 1397 1433 1401
rect 149 1378 157 1382
rect 239 1378 247 1382
rect 780 1376 784 1384
rect 788 1376 792 1384
rect 149 1370 157 1374
rect 239 1370 247 1374
rect 405 1350 413 1354
rect 865 1355 873 1359
rect 1335 1353 1343 1357
rect 1425 1353 1433 1357
rect 865 1347 873 1351
rect 405 1342 413 1346
rect 1335 1345 1343 1349
rect 1425 1345 1433 1349
rect 149 1326 157 1330
rect 239 1326 247 1330
rect 1001 1332 1005 1340
rect 1009 1332 1013 1340
rect 149 1318 157 1322
rect 239 1318 247 1322
rect 48 1306 56 1310
rect 951 1310 959 1314
rect 865 1303 873 1307
rect 951 1302 959 1306
rect 48 1298 56 1302
rect 84 1286 88 1294
rect 92 1286 96 1294
rect 360 1289 368 1293
rect 865 1295 873 1299
rect 360 1281 368 1285
rect 805 1283 813 1287
rect 397 1272 401 1280
rect 405 1272 409 1280
rect 805 1275 813 1279
rect 1331 1279 1339 1283
rect 1421 1279 1429 1283
rect 1331 1271 1339 1275
rect 1421 1271 1429 1275
rect 48 1254 56 1258
rect 48 1246 56 1250
rect 153 1248 161 1252
rect 243 1248 251 1252
rect 865 1260 873 1264
rect 951 1258 959 1262
rect 865 1252 873 1256
rect 951 1250 959 1254
rect -169 1233 -165 1241
rect -161 1233 -157 1241
rect -130 1233 -126 1241
rect -122 1233 -118 1241
rect -90 1233 -86 1241
rect -82 1233 -78 1241
rect -51 1233 -47 1241
rect -43 1233 -39 1241
rect -10 1233 -6 1241
rect -2 1233 2 1241
rect 153 1240 161 1244
rect 243 1240 251 1244
rect 360 1237 368 1241
rect 360 1229 368 1233
rect 1331 1227 1339 1231
rect 1421 1227 1429 1231
rect 1331 1219 1339 1223
rect 1421 1219 1429 1223
rect 865 1208 873 1212
rect 1230 1207 1238 1211
rect 153 1196 161 1200
rect 243 1196 251 1200
rect 865 1200 873 1204
rect 1230 1199 1238 1203
rect 153 1188 161 1192
rect 243 1188 251 1192
rect 320 1183 324 1191
rect 328 1183 332 1191
rect 1266 1187 1270 1195
rect 1274 1187 1278 1195
rect -181 1175 -177 1183
rect -173 1175 -169 1183
rect 405 1162 413 1166
rect 405 1154 413 1158
rect 1230 1155 1238 1159
rect 780 1143 784 1151
rect 788 1143 792 1151
rect 149 1122 157 1126
rect 239 1122 247 1126
rect 1230 1147 1238 1151
rect 1335 1149 1343 1153
rect 1425 1149 1433 1153
rect 1013 1134 1017 1142
rect 1021 1134 1025 1142
rect 1052 1134 1056 1142
rect 1060 1134 1064 1142
rect 1092 1134 1096 1142
rect 1100 1134 1104 1142
rect 1131 1134 1135 1142
rect 1139 1134 1143 1142
rect 1172 1134 1176 1142
rect 1180 1134 1184 1142
rect 1335 1141 1343 1145
rect 1425 1141 1433 1145
rect 149 1114 157 1118
rect 239 1114 247 1118
rect 491 1117 499 1121
rect 865 1122 873 1126
rect 865 1114 873 1118
rect 405 1110 413 1114
rect 491 1109 499 1113
rect 405 1102 413 1106
rect 1335 1097 1343 1101
rect 1425 1097 1433 1101
rect 345 1090 353 1094
rect 345 1082 353 1086
rect 1335 1089 1343 1093
rect 1425 1089 1433 1093
rect 951 1077 959 1081
rect 1001 1076 1005 1084
rect 1009 1076 1013 1084
rect 149 1070 157 1074
rect 239 1070 247 1074
rect 149 1062 157 1066
rect 405 1067 413 1071
rect 865 1070 873 1074
rect 951 1069 959 1073
rect 239 1062 247 1066
rect 491 1065 499 1069
rect 405 1059 413 1063
rect 491 1057 499 1061
rect 865 1062 873 1066
rect 48 1050 56 1054
rect 805 1050 813 1054
rect 48 1042 56 1046
rect 805 1042 813 1046
rect 84 1030 88 1038
rect 92 1030 96 1038
rect 542 1023 546 1031
rect 550 1023 554 1031
rect 580 1023 584 1031
rect 588 1023 592 1031
rect 618 1023 622 1031
rect 626 1023 630 1031
rect 656 1023 660 1031
rect 664 1023 668 1031
rect 725 1024 729 1032
rect 733 1024 737 1032
rect 865 1027 873 1031
rect 951 1025 959 1029
rect 405 1015 413 1019
rect 405 1007 413 1011
rect 865 1019 873 1023
rect 1331 1023 1339 1027
rect 1421 1023 1429 1027
rect 951 1017 959 1021
rect 1331 1015 1339 1019
rect 1421 1015 1429 1019
rect 48 998 56 1002
rect 48 990 56 994
rect 153 992 161 996
rect 243 992 251 996
rect -169 977 -165 985
rect -161 977 -157 985
rect -130 977 -126 985
rect -122 977 -118 985
rect -90 977 -86 985
rect -82 977 -78 985
rect -51 977 -47 985
rect -43 977 -39 985
rect -10 977 -6 985
rect -2 977 2 985
rect 153 984 161 988
rect 243 984 251 988
rect 865 975 873 979
rect 725 967 729 975
rect 733 967 737 975
rect 360 954 368 958
rect 865 967 873 971
rect 1331 971 1339 975
rect 1421 971 1429 975
rect 1331 963 1339 967
rect 1421 963 1429 967
rect 360 946 368 950
rect 153 940 161 944
rect 243 940 251 944
rect 153 932 161 936
rect 243 932 251 936
rect 397 937 401 945
rect 405 937 409 945
rect 1230 951 1238 955
rect 1230 943 1238 947
rect -181 919 -177 927
rect -173 919 -169 927
rect 1266 931 1270 939
rect 1274 931 1278 939
rect 725 910 729 918
rect 733 910 737 918
rect 780 910 784 918
rect 788 910 792 918
rect 360 902 368 906
rect 360 894 368 898
rect 1230 899 1238 903
rect 865 889 873 893
rect 1230 891 1238 895
rect 1335 893 1343 897
rect 1425 893 1433 897
rect 865 881 873 885
rect 149 866 157 870
rect 239 866 247 870
rect 1013 878 1017 886
rect 1021 878 1025 886
rect 1052 878 1056 886
rect 1060 878 1064 886
rect 1092 878 1096 886
rect 1100 878 1104 886
rect 1131 878 1135 886
rect 1139 878 1143 886
rect 1172 878 1176 886
rect 1180 878 1184 886
rect 1335 885 1343 889
rect 1425 885 1433 889
rect 149 858 157 862
rect 239 858 247 862
rect 320 848 324 856
rect 328 848 332 856
rect 725 853 729 861
rect 733 853 737 861
rect 951 844 959 848
rect 1335 841 1343 845
rect 865 837 873 841
rect 1425 841 1433 845
rect 951 836 959 840
rect 405 827 413 831
rect 865 829 873 833
rect 1335 833 1343 837
rect 1425 833 1433 837
rect 405 819 413 823
rect 149 814 157 818
rect 239 814 247 818
rect 805 817 813 821
rect 1001 820 1005 828
rect 1009 820 1013 828
rect 149 806 157 810
rect 239 806 247 810
rect 805 809 813 813
rect 48 794 56 798
rect 48 786 56 790
rect 865 794 873 798
rect 951 792 959 796
rect 865 786 873 790
rect 84 774 88 782
rect 92 774 96 782
rect 491 782 499 786
rect 951 784 959 788
rect 405 775 413 779
rect 491 774 499 778
rect 405 767 413 771
rect 1331 767 1339 771
rect 1421 767 1429 771
rect 345 755 353 759
rect 1331 759 1339 763
rect 1421 759 1429 763
rect 345 747 353 751
rect 48 742 56 746
rect 48 734 56 738
rect 153 736 161 740
rect 865 742 873 746
rect 243 736 251 740
rect -169 721 -165 729
rect -161 721 -157 729
rect -130 721 -126 729
rect -122 721 -118 729
rect -90 721 -86 729
rect -82 721 -78 729
rect -51 721 -47 729
rect -43 721 -39 729
rect -10 721 -6 729
rect -2 721 2 729
rect 153 728 161 732
rect 243 728 251 732
rect 405 732 413 736
rect 491 730 499 734
rect 865 734 873 738
rect 405 724 413 728
rect 491 722 499 726
rect 1331 715 1339 719
rect 1421 715 1429 719
rect 1331 707 1339 711
rect 1421 707 1429 711
rect 1230 695 1238 699
rect 153 684 161 688
rect 243 684 251 688
rect 1230 687 1238 691
rect 153 676 161 680
rect 243 676 251 680
rect 405 680 413 684
rect 780 677 784 685
rect 788 677 792 685
rect -181 663 -177 671
rect -173 663 -169 671
rect 405 672 413 676
rect 1266 675 1270 683
rect 1274 675 1278 683
rect 865 656 873 660
rect 865 648 873 652
rect 1230 643 1238 647
rect 1230 635 1238 639
rect 1335 637 1343 641
rect 1425 637 1433 641
rect 360 619 368 623
rect 1013 622 1017 630
rect 1021 622 1025 630
rect 1052 622 1056 630
rect 1060 622 1064 630
rect 1092 622 1096 630
rect 1100 622 1104 630
rect 1131 622 1135 630
rect 1139 622 1143 630
rect 1172 622 1176 630
rect 1180 622 1184 630
rect 1335 629 1343 633
rect 1425 629 1433 633
rect 149 610 157 614
rect 239 610 247 614
rect 360 611 368 615
rect 951 611 959 615
rect 149 602 157 606
rect 239 602 247 606
rect 397 602 401 610
rect 405 602 409 610
rect 865 604 873 608
rect 951 603 959 607
rect 865 596 873 600
rect 805 584 813 588
rect 1335 585 1343 589
rect 1425 585 1433 589
rect 805 576 813 580
rect 360 567 368 571
rect 1335 577 1343 581
rect 1425 577 1433 581
rect 149 558 157 562
rect 239 558 247 562
rect 360 559 368 563
rect 865 561 873 565
rect 1001 564 1005 572
rect 1009 564 1013 572
rect 951 559 959 563
rect 149 550 157 554
rect 239 550 247 554
rect 865 553 873 557
rect 951 551 959 555
rect 48 538 56 542
rect 48 530 56 534
rect 84 518 88 526
rect 92 518 96 526
rect 320 513 324 521
rect 328 513 332 521
rect 865 509 873 513
rect 1331 511 1339 515
rect 1421 511 1429 515
rect 780 501 784 509
rect 788 501 792 509
rect 405 492 413 496
rect 48 486 56 490
rect 865 501 873 505
rect 1331 503 1339 507
rect 1421 503 1429 507
rect 48 478 56 482
rect 153 480 161 484
rect 405 484 413 488
rect 243 480 251 484
rect -169 465 -165 473
rect -161 465 -157 473
rect -130 465 -126 473
rect -122 465 -118 473
rect -90 465 -86 473
rect -82 465 -78 473
rect -51 465 -47 473
rect -43 465 -39 473
rect -10 465 -6 473
rect -2 465 2 473
rect 153 472 161 476
rect 243 472 251 476
rect 1331 459 1339 463
rect 1421 459 1429 463
rect 491 447 499 451
rect 1331 451 1339 455
rect 1421 451 1429 455
rect 405 440 413 444
rect 491 439 499 443
rect 1230 439 1238 443
rect 153 428 161 432
rect 243 428 251 432
rect 405 432 413 436
rect 1230 431 1238 435
rect 153 420 161 424
rect 243 420 251 424
rect 345 420 353 424
rect 1266 419 1270 427
rect 1274 419 1278 427
rect -181 407 -177 415
rect -173 407 -169 415
rect 345 412 353 416
rect 405 397 413 401
rect 491 395 499 399
rect 405 389 413 393
rect 491 387 499 391
rect 1230 387 1238 391
rect 1230 379 1238 383
rect 1335 381 1343 385
rect 1425 381 1433 385
rect 149 354 157 358
rect 1013 366 1017 374
rect 1021 366 1025 374
rect 1052 366 1056 374
rect 1060 366 1064 374
rect 1092 366 1096 374
rect 1100 366 1104 374
rect 1131 366 1135 374
rect 1139 366 1143 374
rect 1172 366 1176 374
rect 1180 366 1184 374
rect 1335 373 1343 377
rect 1425 373 1433 377
rect 239 354 247 358
rect 149 346 157 350
rect 239 346 247 350
rect 405 345 413 349
rect 405 337 413 341
rect 1335 329 1343 333
rect 1425 329 1433 333
rect 1335 321 1343 325
rect 1425 321 1433 325
rect 1001 308 1005 316
rect 1009 308 1013 316
rect 149 302 157 306
rect 239 302 247 306
rect 149 294 157 298
rect 239 294 247 298
rect 48 282 56 286
rect 360 284 368 288
rect 48 274 56 278
rect 360 276 368 280
rect 84 262 88 270
rect 92 262 96 270
rect 397 267 401 275
rect 405 267 409 275
rect 48 230 56 234
rect 360 232 368 236
rect 48 222 56 226
rect 153 224 161 228
rect 243 224 251 228
rect 360 224 368 228
rect -169 209 -165 217
rect -161 209 -157 217
rect -130 209 -126 217
rect -122 209 -118 217
rect -90 209 -86 217
rect -82 209 -78 217
rect -51 209 -47 217
rect -43 209 -39 217
rect -10 209 -6 217
rect -2 209 2 217
rect 153 216 161 220
rect 243 216 251 220
rect 153 172 161 176
rect 243 172 251 176
rect 153 164 161 168
rect 243 164 251 168
rect -181 151 -177 159
rect -173 151 -169 159
rect 149 98 157 102
rect 239 98 247 102
rect 149 90 157 94
rect 239 90 247 94
rect 149 46 157 50
rect 239 46 247 50
rect 149 38 157 42
rect 239 38 247 42
rect 48 26 56 30
rect 48 18 56 22
rect 84 6 88 14
rect 92 6 96 14
rect 48 -26 56 -22
rect 48 -34 56 -30
rect 153 -32 161 -28
rect 243 -32 251 -28
rect -169 -47 -165 -39
rect -161 -47 -157 -39
rect -130 -47 -126 -39
rect -122 -47 -118 -39
rect -90 -47 -86 -39
rect -82 -47 -78 -39
rect -51 -47 -47 -39
rect -43 -47 -39 -39
rect -10 -47 -6 -39
rect -2 -47 2 -39
rect 153 -40 161 -36
rect 243 -40 251 -36
rect 153 -84 161 -80
rect 243 -84 251 -80
rect 153 -92 161 -88
rect 243 -92 251 -88
rect -181 -105 -177 -97
rect -173 -105 -169 -97
<< polysilicon >>
rect 139 1889 141 1893
rect 229 1889 231 1893
rect 136 1887 149 1889
rect 157 1887 160 1889
rect 226 1887 239 1889
rect 247 1887 250 1889
rect 116 1871 118 1877
rect 206 1871 208 1877
rect 100 1869 103 1871
rect 111 1869 121 1871
rect 190 1869 193 1871
rect 201 1869 211 1871
rect 115 1861 125 1863
rect 133 1861 136 1863
rect 205 1861 215 1863
rect 223 1861 226 1863
rect 119 1852 121 1861
rect 209 1852 211 1861
rect 136 1835 149 1837
rect 157 1835 160 1837
rect 226 1835 239 1837
rect 247 1835 250 1837
rect 139 1831 141 1835
rect 229 1831 231 1835
rect 38 1817 40 1821
rect 35 1815 48 1817
rect 56 1815 59 1817
rect 89 1806 91 1809
rect 15 1799 17 1805
rect -1 1797 2 1799
rect 10 1797 20 1799
rect 14 1789 24 1791
rect 32 1789 35 1791
rect 18 1780 20 1789
rect 89 1790 91 1798
rect 81 1788 91 1790
rect 89 1786 91 1788
rect 89 1775 91 1778
rect 35 1763 48 1765
rect 56 1763 59 1765
rect 38 1759 40 1763
rect -164 1753 -162 1756
rect -125 1753 -123 1756
rect -85 1753 -83 1756
rect -46 1753 -44 1756
rect -5 1753 -3 1756
rect 143 1759 145 1763
rect 233 1759 235 1763
rect 140 1757 153 1759
rect 161 1757 164 1759
rect 230 1757 243 1759
rect 251 1757 254 1759
rect -164 1737 -162 1745
rect -172 1735 -162 1737
rect -164 1733 -162 1735
rect -125 1737 -123 1745
rect -133 1735 -123 1737
rect -125 1733 -123 1735
rect -85 1737 -83 1745
rect -93 1735 -83 1737
rect -85 1733 -83 1735
rect -46 1737 -44 1745
rect -54 1735 -44 1737
rect -46 1733 -44 1735
rect -5 1737 -3 1745
rect 120 1741 122 1747
rect 210 1741 212 1747
rect 104 1739 107 1741
rect 115 1739 125 1741
rect 194 1739 197 1741
rect 205 1739 215 1741
rect -13 1735 -3 1737
rect -5 1733 -3 1735
rect 119 1731 129 1733
rect 137 1731 140 1733
rect 209 1731 219 1733
rect 227 1731 230 1733
rect -164 1722 -162 1725
rect -125 1722 -123 1725
rect -85 1722 -83 1725
rect -46 1722 -44 1725
rect -5 1722 -3 1725
rect 123 1722 125 1731
rect 213 1722 215 1731
rect 140 1705 153 1707
rect 161 1705 164 1707
rect 230 1705 243 1707
rect 251 1705 254 1707
rect 143 1701 145 1705
rect -176 1695 -174 1698
rect 233 1701 235 1705
rect -176 1679 -174 1687
rect -184 1677 -174 1679
rect -176 1675 -174 1677
rect -176 1664 -174 1667
rect 139 1633 141 1637
rect 229 1633 231 1637
rect 136 1631 149 1633
rect 157 1631 160 1633
rect 226 1631 239 1633
rect 247 1631 250 1633
rect 116 1615 118 1621
rect 206 1615 208 1621
rect 100 1613 103 1615
rect 111 1613 121 1615
rect 190 1613 193 1615
rect 201 1613 211 1615
rect 115 1605 125 1607
rect 133 1605 136 1607
rect 205 1605 215 1607
rect 223 1605 226 1607
rect 119 1596 121 1605
rect 209 1596 211 1605
rect 136 1579 149 1581
rect 157 1579 160 1581
rect 226 1579 239 1581
rect 247 1579 250 1581
rect 139 1575 141 1579
rect 229 1575 231 1579
rect 38 1561 40 1565
rect 35 1559 48 1561
rect 56 1559 59 1561
rect 89 1550 91 1553
rect 15 1543 17 1549
rect -1 1541 2 1543
rect 10 1541 20 1543
rect 14 1533 24 1535
rect 32 1533 35 1535
rect 18 1524 20 1533
rect 89 1534 91 1542
rect 1321 1534 1323 1538
rect 1411 1534 1413 1538
rect 81 1532 91 1534
rect 1318 1532 1331 1534
rect 1339 1532 1342 1534
rect 1408 1532 1421 1534
rect 1429 1532 1432 1534
rect 89 1530 91 1532
rect 325 1526 327 1529
rect 89 1519 91 1522
rect 35 1507 48 1509
rect 56 1507 59 1509
rect 38 1503 40 1507
rect -164 1497 -162 1500
rect -125 1497 -123 1500
rect -85 1497 -83 1500
rect -46 1497 -44 1500
rect -5 1497 -3 1500
rect 143 1503 145 1507
rect 233 1503 235 1507
rect 325 1510 327 1518
rect 1298 1516 1300 1522
rect 1388 1516 1390 1522
rect 1282 1514 1285 1516
rect 1293 1514 1303 1516
rect 1372 1514 1375 1516
rect 1383 1514 1393 1516
rect 317 1508 327 1510
rect 325 1506 327 1508
rect 1297 1506 1307 1508
rect 1315 1506 1318 1508
rect 1387 1506 1397 1508
rect 1405 1506 1408 1508
rect 140 1501 153 1503
rect 161 1501 164 1503
rect 230 1501 243 1503
rect 251 1501 254 1503
rect 325 1495 327 1498
rect 395 1496 397 1500
rect 1301 1497 1303 1506
rect 1391 1497 1393 1506
rect 392 1494 405 1496
rect 413 1494 416 1496
rect -164 1481 -162 1489
rect -172 1479 -162 1481
rect -164 1477 -162 1479
rect -125 1481 -123 1489
rect -133 1479 -123 1481
rect -125 1477 -123 1479
rect -85 1481 -83 1489
rect -93 1479 -83 1481
rect -85 1477 -83 1479
rect -46 1481 -44 1489
rect -54 1479 -44 1481
rect -46 1477 -44 1479
rect -5 1481 -3 1489
rect 120 1485 122 1491
rect 210 1485 212 1491
rect 104 1483 107 1485
rect 115 1483 125 1485
rect 194 1483 197 1485
rect 205 1483 215 1485
rect -13 1479 -3 1481
rect -5 1477 -3 1479
rect 372 1478 374 1484
rect 1318 1480 1331 1482
rect 1339 1480 1342 1482
rect 1408 1480 1421 1482
rect 1429 1480 1432 1482
rect 119 1475 129 1477
rect 137 1475 140 1477
rect 209 1475 219 1477
rect 227 1475 230 1477
rect 356 1476 359 1478
rect 367 1476 377 1478
rect 1321 1476 1323 1480
rect -164 1466 -162 1469
rect -125 1466 -123 1469
rect -85 1466 -83 1469
rect -46 1466 -44 1469
rect -5 1466 -3 1469
rect 123 1466 125 1475
rect 213 1466 215 1475
rect 1411 1476 1413 1480
rect 371 1468 381 1470
rect 389 1468 392 1470
rect 375 1459 377 1468
rect 1220 1462 1222 1466
rect 1217 1460 1230 1462
rect 1238 1460 1241 1462
rect 481 1451 483 1455
rect 140 1449 153 1451
rect 161 1449 164 1451
rect 230 1449 243 1451
rect 251 1449 254 1451
rect 478 1449 491 1451
rect 499 1449 502 1451
rect 1271 1451 1273 1454
rect 143 1445 145 1449
rect -176 1439 -174 1442
rect 233 1445 235 1449
rect 1197 1444 1199 1450
rect 392 1442 405 1444
rect 413 1442 416 1444
rect 395 1438 397 1442
rect 1181 1442 1184 1444
rect 1192 1442 1202 1444
rect 458 1433 460 1439
rect 1196 1434 1206 1436
rect 1214 1434 1217 1436
rect -176 1423 -174 1431
rect 335 1424 337 1432
rect 442 1431 445 1433
rect 453 1431 463 1433
rect 1200 1425 1202 1434
rect 1271 1435 1273 1443
rect 1263 1433 1273 1435
rect 1271 1431 1273 1433
rect -184 1421 -174 1423
rect 322 1422 325 1424
rect 333 1422 345 1424
rect 353 1422 356 1424
rect 457 1423 467 1425
rect 475 1423 478 1425
rect -176 1419 -174 1421
rect 461 1414 463 1423
rect 1271 1420 1273 1423
rect -176 1408 -174 1411
rect 1217 1408 1230 1410
rect 1238 1408 1241 1410
rect 395 1401 397 1405
rect 1220 1404 1222 1408
rect 392 1399 405 1401
rect 413 1399 416 1401
rect 478 1397 491 1399
rect 499 1397 502 1399
rect 1018 1398 1020 1401
rect 1057 1398 1059 1401
rect 1097 1398 1099 1401
rect 1136 1398 1138 1401
rect 1177 1398 1179 1401
rect 1325 1404 1327 1408
rect 1415 1404 1417 1408
rect 1322 1402 1335 1404
rect 1343 1402 1346 1404
rect 1412 1402 1425 1404
rect 1433 1402 1436 1404
rect 481 1393 483 1397
rect 139 1377 141 1381
rect 372 1383 374 1389
rect 785 1384 787 1387
rect 229 1377 231 1381
rect 356 1381 359 1383
rect 367 1381 377 1383
rect 136 1375 149 1377
rect 157 1375 160 1377
rect 226 1375 239 1377
rect 247 1375 250 1377
rect 1018 1382 1020 1390
rect 1010 1380 1020 1382
rect 1018 1378 1020 1380
rect 1057 1382 1059 1390
rect 1049 1380 1059 1382
rect 1057 1378 1059 1380
rect 1097 1382 1099 1390
rect 1089 1380 1099 1382
rect 1097 1378 1099 1380
rect 1136 1382 1138 1390
rect 1128 1380 1138 1382
rect 1136 1378 1138 1380
rect 1177 1382 1179 1390
rect 1302 1386 1304 1392
rect 1392 1386 1394 1392
rect 1286 1384 1289 1386
rect 1297 1384 1307 1386
rect 1376 1384 1379 1386
rect 1387 1384 1397 1386
rect 1169 1380 1179 1382
rect 1177 1378 1179 1380
rect 371 1373 381 1375
rect 389 1373 392 1375
rect 116 1359 118 1365
rect 206 1359 208 1365
rect 375 1364 377 1373
rect 785 1368 787 1376
rect 1301 1376 1311 1378
rect 1319 1376 1322 1378
rect 1391 1376 1401 1378
rect 1409 1376 1412 1378
rect 777 1366 787 1368
rect 1018 1367 1020 1370
rect 1057 1367 1059 1370
rect 1097 1367 1099 1370
rect 1136 1367 1138 1370
rect 1177 1367 1179 1370
rect 1305 1367 1307 1376
rect 1395 1367 1397 1376
rect 785 1364 787 1366
rect 100 1357 103 1359
rect 111 1357 121 1359
rect 190 1357 193 1359
rect 201 1357 211 1359
rect 115 1349 125 1351
rect 133 1349 136 1351
rect 205 1349 215 1351
rect 223 1349 226 1351
rect 785 1353 787 1356
rect 855 1354 857 1358
rect 852 1352 865 1354
rect 873 1352 876 1354
rect 119 1340 121 1349
rect 209 1340 211 1349
rect 392 1347 405 1349
rect 413 1347 416 1349
rect 1322 1350 1335 1352
rect 1343 1350 1346 1352
rect 1412 1350 1425 1352
rect 1433 1350 1436 1352
rect 395 1343 397 1347
rect 1325 1346 1327 1350
rect 832 1336 834 1342
rect 1006 1340 1008 1343
rect 1415 1346 1417 1350
rect 816 1334 819 1336
rect 827 1334 837 1336
rect 831 1326 841 1328
rect 849 1326 852 1328
rect 136 1323 149 1325
rect 157 1323 160 1325
rect 226 1323 239 1325
rect 247 1323 250 1325
rect 139 1319 141 1323
rect 229 1319 231 1323
rect 835 1317 837 1326
rect 1006 1324 1008 1332
rect 998 1322 1008 1324
rect 1006 1320 1008 1322
rect 38 1305 40 1309
rect 941 1309 943 1313
rect 1006 1309 1008 1312
rect 938 1307 951 1309
rect 959 1307 962 1309
rect 35 1303 48 1305
rect 56 1303 59 1305
rect 852 1300 865 1302
rect 873 1300 876 1302
rect 89 1294 91 1297
rect 855 1296 857 1300
rect 15 1287 17 1293
rect -1 1285 2 1287
rect 10 1285 20 1287
rect 350 1288 352 1292
rect 918 1291 920 1297
rect 347 1286 360 1288
rect 368 1286 371 1288
rect 14 1277 24 1279
rect 32 1277 35 1279
rect 18 1268 20 1277
rect 89 1278 91 1286
rect 402 1280 404 1283
rect 795 1282 797 1290
rect 902 1289 905 1291
rect 913 1289 923 1291
rect 782 1280 785 1282
rect 793 1280 805 1282
rect 813 1280 816 1282
rect 917 1281 927 1283
rect 935 1281 938 1283
rect 81 1276 91 1278
rect 89 1274 91 1276
rect 327 1270 329 1276
rect 921 1272 923 1281
rect 1321 1278 1323 1282
rect 1411 1278 1413 1282
rect 1318 1276 1331 1278
rect 1339 1276 1342 1278
rect 1408 1276 1421 1278
rect 1429 1276 1432 1278
rect 311 1268 314 1270
rect 322 1268 332 1270
rect 89 1263 91 1266
rect 326 1260 336 1262
rect 344 1260 347 1262
rect 402 1264 404 1272
rect 394 1262 404 1264
rect 402 1260 404 1262
rect 35 1251 48 1253
rect 56 1251 59 1253
rect 38 1247 40 1251
rect -164 1241 -162 1244
rect -125 1241 -123 1244
rect -85 1241 -83 1244
rect -46 1241 -44 1244
rect -5 1241 -3 1244
rect 143 1247 145 1251
rect 233 1247 235 1251
rect 330 1251 332 1260
rect 855 1259 857 1263
rect 852 1257 865 1259
rect 873 1257 876 1259
rect 1298 1260 1300 1266
rect 1388 1260 1390 1266
rect 1282 1258 1285 1260
rect 1293 1258 1303 1260
rect 1372 1258 1375 1260
rect 1383 1258 1393 1260
rect 938 1255 951 1257
rect 959 1255 962 1257
rect 402 1249 404 1252
rect 941 1251 943 1255
rect 1297 1250 1307 1252
rect 1315 1250 1318 1252
rect 1387 1250 1397 1252
rect 1405 1250 1408 1252
rect 140 1245 153 1247
rect 161 1245 164 1247
rect 230 1245 243 1247
rect 251 1245 254 1247
rect 832 1241 834 1247
rect 1301 1241 1303 1250
rect 1391 1241 1393 1250
rect 816 1239 819 1241
rect 827 1239 837 1241
rect -164 1225 -162 1233
rect -172 1223 -162 1225
rect -164 1221 -162 1223
rect -125 1225 -123 1233
rect -133 1223 -123 1225
rect -125 1221 -123 1223
rect -85 1225 -83 1233
rect -93 1223 -83 1225
rect -85 1221 -83 1223
rect -46 1225 -44 1233
rect -54 1223 -44 1225
rect -46 1221 -44 1223
rect -5 1225 -3 1233
rect 120 1229 122 1235
rect 210 1229 212 1235
rect 347 1234 360 1236
rect 368 1234 371 1236
rect 350 1230 352 1234
rect 104 1227 107 1229
rect 115 1227 125 1229
rect 194 1227 197 1229
rect 205 1227 215 1229
rect -13 1223 -3 1225
rect -5 1221 -3 1223
rect 831 1231 841 1233
rect 849 1231 852 1233
rect 835 1222 837 1231
rect 1318 1224 1331 1226
rect 1339 1224 1342 1226
rect 1408 1224 1421 1226
rect 1429 1224 1432 1226
rect 119 1219 129 1221
rect 137 1219 140 1221
rect 209 1219 219 1221
rect 227 1219 230 1221
rect -164 1210 -162 1213
rect -125 1210 -123 1213
rect -85 1210 -83 1213
rect -46 1210 -44 1213
rect -5 1210 -3 1213
rect 123 1210 125 1219
rect 213 1210 215 1219
rect 1321 1220 1323 1224
rect 1411 1220 1413 1224
rect 852 1205 865 1207
rect 873 1205 876 1207
rect 1220 1206 1222 1210
rect 855 1201 857 1205
rect 1217 1204 1230 1206
rect 1238 1204 1241 1206
rect 140 1193 153 1195
rect 161 1193 164 1195
rect 230 1193 243 1195
rect 251 1193 254 1195
rect 1271 1195 1273 1198
rect 143 1189 145 1193
rect -176 1183 -174 1186
rect 233 1189 235 1193
rect 325 1191 327 1194
rect 1197 1188 1199 1194
rect 1181 1186 1184 1188
rect 1192 1186 1202 1188
rect -176 1167 -174 1175
rect 325 1175 327 1183
rect 1196 1178 1206 1180
rect 1214 1178 1217 1180
rect 317 1173 327 1175
rect 325 1171 327 1173
rect -184 1165 -174 1167
rect -176 1163 -174 1165
rect 1200 1169 1202 1178
rect 1271 1179 1273 1187
rect 1263 1177 1273 1179
rect 1271 1175 1273 1177
rect 325 1160 327 1163
rect 395 1161 397 1165
rect 1271 1164 1273 1167
rect 392 1159 405 1161
rect 413 1159 416 1161
rect -176 1152 -174 1155
rect 785 1151 787 1154
rect 1217 1152 1230 1154
rect 1238 1152 1241 1154
rect 372 1143 374 1149
rect 1220 1148 1222 1152
rect 356 1141 359 1143
rect 367 1141 377 1143
rect 371 1133 381 1135
rect 389 1133 392 1135
rect 139 1121 141 1125
rect 229 1121 231 1125
rect 375 1124 377 1133
rect 785 1135 787 1143
rect 1018 1142 1020 1145
rect 1057 1142 1059 1145
rect 1097 1142 1099 1145
rect 1136 1142 1138 1145
rect 1177 1142 1179 1145
rect 1325 1148 1327 1152
rect 1415 1148 1417 1152
rect 1322 1146 1335 1148
rect 1343 1146 1346 1148
rect 1412 1146 1425 1148
rect 1433 1146 1436 1148
rect 777 1133 787 1135
rect 785 1131 787 1133
rect 136 1119 149 1121
rect 157 1119 160 1121
rect 226 1119 239 1121
rect 247 1119 250 1121
rect 481 1116 483 1120
rect 785 1120 787 1123
rect 855 1121 857 1125
rect 1018 1126 1020 1134
rect 1010 1124 1020 1126
rect 1018 1122 1020 1124
rect 1057 1126 1059 1134
rect 1049 1124 1059 1126
rect 1057 1122 1059 1124
rect 1097 1126 1099 1134
rect 1089 1124 1099 1126
rect 1097 1122 1099 1124
rect 1136 1126 1138 1134
rect 1128 1124 1138 1126
rect 1136 1122 1138 1124
rect 1177 1126 1179 1134
rect 1302 1130 1304 1136
rect 1392 1130 1394 1136
rect 1286 1128 1289 1130
rect 1297 1128 1307 1130
rect 1376 1128 1379 1130
rect 1387 1128 1397 1130
rect 1169 1124 1179 1126
rect 1177 1122 1179 1124
rect 852 1119 865 1121
rect 873 1119 876 1121
rect 478 1114 491 1116
rect 499 1114 502 1116
rect 1301 1120 1311 1122
rect 1319 1120 1322 1122
rect 1391 1120 1401 1122
rect 1409 1120 1412 1122
rect 1018 1111 1020 1114
rect 1057 1111 1059 1114
rect 1097 1111 1099 1114
rect 1136 1111 1138 1114
rect 1177 1111 1179 1114
rect 1305 1111 1307 1120
rect 1395 1111 1397 1120
rect 116 1103 118 1109
rect 206 1103 208 1109
rect 392 1107 405 1109
rect 413 1107 416 1109
rect 395 1103 397 1107
rect 100 1101 103 1103
rect 111 1101 121 1103
rect 190 1101 193 1103
rect 201 1101 211 1103
rect 458 1098 460 1104
rect 832 1103 834 1109
rect 816 1101 819 1103
rect 827 1101 837 1103
rect 115 1093 125 1095
rect 133 1093 136 1095
rect 205 1093 215 1095
rect 223 1093 226 1095
rect 119 1084 121 1093
rect 209 1084 211 1093
rect 335 1089 337 1097
rect 442 1096 445 1098
rect 453 1096 463 1098
rect 831 1093 841 1095
rect 849 1093 852 1095
rect 1322 1094 1335 1096
rect 1343 1094 1346 1096
rect 1412 1094 1425 1096
rect 1433 1094 1436 1096
rect 322 1087 325 1089
rect 333 1087 345 1089
rect 353 1087 356 1089
rect 457 1088 467 1090
rect 475 1088 478 1090
rect 461 1079 463 1088
rect 835 1084 837 1093
rect 1325 1090 1327 1094
rect 1006 1084 1008 1087
rect 1415 1090 1417 1094
rect 941 1076 943 1080
rect 938 1074 951 1076
rect 959 1074 962 1076
rect 136 1067 149 1069
rect 157 1067 160 1069
rect 226 1067 239 1069
rect 247 1067 250 1069
rect 139 1063 141 1067
rect 229 1063 231 1067
rect 395 1066 397 1070
rect 392 1064 405 1066
rect 413 1064 416 1066
rect 852 1067 865 1069
rect 873 1067 876 1069
rect 478 1062 491 1064
rect 499 1062 502 1064
rect 855 1063 857 1067
rect 481 1058 483 1062
rect 1006 1068 1008 1076
rect 998 1066 1008 1068
rect 1006 1064 1008 1066
rect 918 1058 920 1064
rect 38 1049 40 1053
rect 35 1047 48 1049
rect 56 1047 59 1049
rect 372 1048 374 1054
rect 795 1049 797 1057
rect 902 1056 905 1058
rect 913 1056 923 1058
rect 1006 1053 1008 1056
rect 356 1046 359 1048
rect 367 1046 377 1048
rect 782 1047 785 1049
rect 793 1047 805 1049
rect 813 1047 816 1049
rect 917 1048 927 1050
rect 935 1048 938 1050
rect 89 1038 91 1041
rect 371 1038 381 1040
rect 389 1038 392 1040
rect 921 1039 923 1048
rect 15 1031 17 1037
rect -1 1029 2 1031
rect 10 1029 20 1031
rect 14 1021 24 1023
rect 32 1021 35 1023
rect 18 1012 20 1021
rect 89 1022 91 1030
rect 375 1029 377 1038
rect 547 1031 549 1034
rect 585 1031 587 1034
rect 623 1031 625 1034
rect 661 1031 663 1034
rect 730 1032 732 1035
rect 855 1026 857 1030
rect 852 1024 865 1026
rect 873 1024 876 1026
rect 81 1020 91 1022
rect 89 1018 91 1020
rect 392 1012 405 1014
rect 413 1012 416 1014
rect 547 1015 549 1023
rect 543 1013 549 1015
rect 89 1007 91 1010
rect 395 1008 397 1012
rect 547 1010 549 1013
rect 585 1015 587 1023
rect 581 1013 587 1015
rect 585 1010 587 1013
rect 623 1015 625 1023
rect 619 1013 625 1015
rect 623 1010 625 1013
rect 661 1015 663 1023
rect 657 1013 663 1015
rect 730 1016 732 1024
rect 938 1022 951 1024
rect 959 1022 962 1024
rect 1321 1022 1323 1026
rect 1411 1022 1413 1026
rect 941 1018 943 1022
rect 722 1014 732 1016
rect 1318 1020 1331 1022
rect 1339 1020 1342 1022
rect 1408 1020 1421 1022
rect 1429 1020 1432 1022
rect 661 1010 663 1013
rect 730 1012 732 1014
rect 832 1008 834 1014
rect 816 1006 819 1008
rect 827 1006 837 1008
rect 730 1001 732 1004
rect 1298 1004 1300 1010
rect 1388 1004 1390 1010
rect 1282 1002 1285 1004
rect 1293 1002 1303 1004
rect 1372 1002 1375 1004
rect 1383 1002 1393 1004
rect 35 995 48 997
rect 56 995 59 997
rect 38 991 40 995
rect -164 985 -162 988
rect -125 985 -123 988
rect -85 985 -83 988
rect -46 985 -44 988
rect -5 985 -3 988
rect 143 991 145 995
rect 831 998 841 1000
rect 849 998 852 1000
rect 233 991 235 995
rect 661 991 663 994
rect 691 992 693 995
rect 140 989 153 991
rect 161 989 164 991
rect 230 989 243 991
rect 251 989 254 991
rect 835 989 837 998
rect 1297 994 1307 996
rect 1315 994 1318 996
rect 1387 994 1397 996
rect 1405 994 1408 996
rect 1301 985 1303 994
rect 1391 985 1393 994
rect 661 979 663 983
rect 691 980 693 984
rect -164 969 -162 977
rect -172 967 -162 969
rect -164 965 -162 967
rect -125 969 -123 977
rect -133 967 -123 969
rect -125 965 -123 967
rect -85 969 -83 977
rect -93 967 -83 969
rect -85 965 -83 967
rect -46 969 -44 977
rect -54 967 -44 969
rect -46 965 -44 967
rect -5 969 -3 977
rect 120 973 122 979
rect 210 973 212 979
rect 661 977 672 979
rect 661 973 663 977
rect 691 978 702 980
rect 691 974 693 978
rect 730 975 732 978
rect 104 971 107 973
rect 115 971 125 973
rect 194 971 197 973
rect 205 971 215 973
rect -13 967 -3 969
rect -5 965 -3 967
rect 653 968 655 971
rect 647 966 655 968
rect 852 972 865 974
rect 873 972 876 974
rect 855 968 857 972
rect 119 963 129 965
rect 137 963 140 965
rect 209 963 219 965
rect 227 963 230 965
rect -164 954 -162 957
rect -125 954 -123 957
rect -85 954 -83 957
rect -46 954 -44 957
rect -5 954 -3 957
rect 123 954 125 963
rect 213 954 215 963
rect 653 961 655 966
rect 350 953 352 957
rect 730 959 732 967
rect 1318 968 1331 970
rect 1339 968 1342 970
rect 1408 968 1421 970
rect 1429 968 1432 970
rect 1321 964 1323 968
rect 1411 964 1413 968
rect 722 957 732 959
rect 730 955 732 957
rect 347 951 360 953
rect 368 951 371 953
rect 623 950 625 953
rect 653 950 655 953
rect 402 945 404 948
rect 140 937 153 939
rect 161 937 164 939
rect 230 937 243 939
rect 251 937 254 939
rect 143 933 145 937
rect -176 927 -174 930
rect 233 933 235 937
rect 327 935 329 941
rect 1220 950 1222 954
rect 1217 948 1230 950
rect 1238 948 1241 950
rect 730 944 732 947
rect 623 938 625 942
rect 311 933 314 935
rect 322 933 332 935
rect 326 925 336 927
rect 344 925 347 927
rect 402 929 404 937
rect 623 936 634 938
rect 623 932 625 936
rect 1271 939 1273 942
rect 1197 932 1199 938
rect 1181 930 1184 932
rect 1192 930 1202 932
rect 394 927 404 929
rect 402 925 404 927
rect -176 911 -174 919
rect 330 916 332 925
rect 615 927 617 930
rect 609 925 617 927
rect 615 920 617 925
rect 1196 922 1206 924
rect 1214 922 1217 924
rect 402 914 404 917
rect 730 918 732 921
rect 785 918 787 921
rect -184 909 -174 911
rect 585 909 587 912
rect 615 909 617 912
rect 1200 913 1202 922
rect 1271 923 1273 931
rect 1263 921 1273 923
rect 1271 919 1273 921
rect -176 907 -174 909
rect 347 899 360 901
rect 368 899 371 901
rect -176 896 -174 899
rect 350 895 352 899
rect 585 897 587 901
rect 730 902 732 910
rect 722 900 732 902
rect 730 898 732 900
rect 785 902 787 910
rect 1271 908 1273 911
rect 777 900 787 902
rect 785 898 787 900
rect 585 895 596 897
rect 585 891 587 895
rect 1217 896 1230 898
rect 1238 896 1241 898
rect 577 886 579 889
rect 730 887 732 890
rect 785 887 787 890
rect 855 888 857 892
rect 1220 892 1222 896
rect 852 886 865 888
rect 873 886 876 888
rect 1018 886 1020 889
rect 1057 886 1059 889
rect 1097 886 1099 889
rect 1136 886 1138 889
rect 1177 886 1179 889
rect 1325 892 1327 896
rect 1415 892 1417 896
rect 1322 890 1335 892
rect 1343 890 1346 892
rect 1412 890 1425 892
rect 1433 890 1436 892
rect 571 884 579 886
rect 577 879 579 884
rect 139 865 141 869
rect 547 875 549 878
rect 541 873 549 875
rect 229 865 231 869
rect 547 868 549 873
rect 577 868 579 871
rect 832 870 834 876
rect 816 868 819 870
rect 827 868 837 870
rect 136 863 149 865
rect 157 863 160 865
rect 226 863 239 865
rect 247 863 250 865
rect 1018 870 1020 878
rect 1010 868 1020 870
rect 730 861 732 864
rect 1018 866 1020 868
rect 1057 870 1059 878
rect 1049 868 1059 870
rect 1057 866 1059 868
rect 1097 870 1099 878
rect 1089 868 1099 870
rect 1097 866 1099 868
rect 1136 870 1138 878
rect 1128 868 1138 870
rect 1136 866 1138 868
rect 1177 870 1179 878
rect 1302 874 1304 880
rect 1392 874 1394 880
rect 1286 872 1289 874
rect 1297 872 1307 874
rect 1376 872 1379 874
rect 1387 872 1397 874
rect 1169 868 1179 870
rect 1177 866 1179 868
rect 325 856 327 859
rect 547 857 549 860
rect 116 847 118 853
rect 206 847 208 853
rect 831 860 841 862
rect 849 860 852 862
rect 100 845 103 847
rect 111 845 121 847
rect 190 845 193 847
rect 201 845 211 847
rect 115 837 125 839
rect 133 837 136 839
rect 205 837 215 839
rect 223 837 226 839
rect 325 840 327 848
rect 539 846 541 849
rect 533 844 541 846
rect 317 838 327 840
rect 539 839 541 844
rect 730 845 732 853
rect 835 851 837 860
rect 1301 864 1311 866
rect 1319 864 1322 866
rect 1391 864 1401 866
rect 1409 864 1412 866
rect 1018 855 1020 858
rect 1057 855 1059 858
rect 1097 855 1099 858
rect 1136 855 1138 858
rect 1177 855 1179 858
rect 1305 855 1307 864
rect 1395 855 1397 864
rect 722 843 732 845
rect 941 843 943 847
rect 730 841 732 843
rect 938 841 951 843
rect 959 841 962 843
rect 119 828 121 837
rect 209 828 211 837
rect 325 836 327 838
rect 1322 838 1335 840
rect 1343 838 1346 840
rect 1412 838 1425 840
rect 1433 838 1436 840
rect 852 834 865 836
rect 873 834 876 836
rect 325 825 327 828
rect 395 826 397 830
rect 539 828 541 831
rect 730 830 732 833
rect 855 830 857 834
rect 392 824 405 826
rect 413 824 416 826
rect 1325 834 1327 838
rect 918 825 920 831
rect 1006 828 1008 831
rect 1415 834 1417 838
rect 531 817 533 820
rect 525 815 533 817
rect 795 816 797 824
rect 902 823 905 825
rect 913 823 923 825
rect 136 811 149 813
rect 157 811 160 813
rect 226 811 239 813
rect 247 811 250 813
rect 139 807 141 811
rect 229 807 231 811
rect 372 808 374 814
rect 531 810 533 815
rect 782 814 785 816
rect 793 814 805 816
rect 813 814 816 816
rect 917 815 927 817
rect 935 815 938 817
rect 356 806 359 808
rect 367 806 377 808
rect 921 806 923 815
rect 1006 812 1008 820
rect 998 810 1008 812
rect 1006 808 1008 810
rect 371 798 381 800
rect 389 798 392 800
rect 531 799 533 802
rect 38 793 40 797
rect 35 791 48 793
rect 56 791 59 793
rect 375 789 377 798
rect 855 793 857 797
rect 1006 797 1008 800
rect 852 791 865 793
rect 873 791 876 793
rect 938 789 951 791
rect 959 789 962 791
rect 89 782 91 785
rect 15 775 17 781
rect -1 773 2 775
rect 10 773 20 775
rect 481 781 483 785
rect 941 785 943 789
rect 478 779 491 781
rect 499 779 502 781
rect 832 775 834 781
rect 14 765 24 767
rect 32 765 35 767
rect 18 756 20 765
rect 89 766 91 774
rect 392 772 405 774
rect 413 772 416 774
rect 816 773 819 775
rect 827 773 837 775
rect 395 768 397 772
rect 81 764 91 766
rect 89 762 91 764
rect 458 763 460 769
rect 831 765 841 767
rect 849 765 852 767
rect 1321 766 1323 770
rect 1411 766 1413 770
rect 335 754 337 762
rect 442 761 445 763
rect 453 761 463 763
rect 835 756 837 765
rect 1318 764 1331 766
rect 1339 764 1342 766
rect 1408 764 1421 766
rect 1429 764 1432 766
rect 89 751 91 754
rect 322 752 325 754
rect 333 752 345 754
rect 353 752 356 754
rect 457 753 467 755
rect 475 753 478 755
rect 461 744 463 753
rect 1298 748 1300 754
rect 1388 748 1390 754
rect 1282 746 1285 748
rect 1293 746 1303 748
rect 1372 746 1375 748
rect 1383 746 1393 748
rect 35 739 48 741
rect 56 739 59 741
rect 38 735 40 739
rect -164 729 -162 732
rect -125 729 -123 732
rect -85 729 -83 732
rect -46 729 -44 732
rect -5 729 -3 732
rect 143 735 145 739
rect 233 735 235 739
rect 852 739 865 741
rect 873 739 876 741
rect 140 733 153 735
rect 161 733 164 735
rect 230 733 243 735
rect 251 733 254 735
rect 395 731 397 735
rect 855 735 857 739
rect 1297 738 1307 740
rect 1315 738 1318 740
rect 1387 738 1397 740
rect 1405 738 1408 740
rect 392 729 405 731
rect 413 729 416 731
rect 1301 729 1303 738
rect 1391 729 1393 738
rect 478 727 491 729
rect 499 727 502 729
rect 481 723 483 727
rect -164 713 -162 721
rect -172 711 -162 713
rect -164 709 -162 711
rect -125 713 -123 721
rect -133 711 -123 713
rect -125 709 -123 711
rect -85 713 -83 721
rect -93 711 -83 713
rect -85 709 -83 711
rect -46 713 -44 721
rect -54 711 -44 713
rect -46 709 -44 711
rect -5 713 -3 721
rect 120 717 122 723
rect 210 717 212 723
rect 104 715 107 717
rect 115 715 125 717
rect 194 715 197 717
rect 205 715 215 717
rect -13 711 -3 713
rect -5 709 -3 711
rect 372 713 374 719
rect 356 711 359 713
rect 367 711 377 713
rect 1318 712 1331 714
rect 1339 712 1342 714
rect 1408 712 1421 714
rect 1429 712 1432 714
rect 119 707 129 709
rect 137 707 140 709
rect 209 707 219 709
rect 227 707 230 709
rect -164 698 -162 701
rect -125 698 -123 701
rect -85 698 -83 701
rect -46 698 -44 701
rect -5 698 -3 701
rect 123 698 125 707
rect 213 698 215 707
rect 1321 708 1323 712
rect 371 703 381 705
rect 389 703 392 705
rect 1411 708 1413 712
rect 375 694 377 703
rect 1220 694 1222 698
rect 1217 692 1230 694
rect 1238 692 1241 694
rect 785 685 787 688
rect 140 681 153 683
rect 161 681 164 683
rect 230 681 243 683
rect 251 681 254 683
rect 143 677 145 681
rect -176 671 -174 674
rect 233 677 235 681
rect 392 677 405 679
rect 413 677 416 679
rect 1271 683 1273 686
rect 395 673 397 677
rect 785 669 787 677
rect 1197 676 1199 682
rect 1181 674 1184 676
rect 1192 674 1202 676
rect 777 667 787 669
rect 785 665 787 667
rect 1196 666 1206 668
rect 1214 666 1217 668
rect -176 655 -174 663
rect -184 653 -174 655
rect 785 654 787 657
rect 855 655 857 659
rect 1200 657 1202 666
rect 1271 667 1273 675
rect 1263 665 1273 667
rect 1271 663 1273 665
rect 852 653 865 655
rect 873 653 876 655
rect -176 651 -174 653
rect 1271 652 1273 655
rect -176 640 -174 643
rect 832 637 834 643
rect 1217 640 1230 642
rect 1238 640 1241 642
rect 816 635 819 637
rect 827 635 837 637
rect 1220 636 1222 640
rect 1018 630 1020 633
rect 1057 630 1059 633
rect 1097 630 1099 633
rect 1136 630 1138 633
rect 1177 630 1179 633
rect 1325 636 1327 640
rect 1415 636 1417 640
rect 1322 634 1335 636
rect 1343 634 1346 636
rect 1412 634 1425 636
rect 1433 634 1436 636
rect 831 627 841 629
rect 849 627 852 629
rect 350 618 352 622
rect 835 618 837 627
rect 139 609 141 613
rect 347 616 360 618
rect 368 616 371 618
rect 229 609 231 613
rect 402 610 404 613
rect 941 610 943 614
rect 1018 614 1020 622
rect 1010 612 1020 614
rect 1018 610 1020 612
rect 1057 614 1059 622
rect 1049 612 1059 614
rect 1057 610 1059 612
rect 1097 614 1099 622
rect 1089 612 1099 614
rect 1097 610 1099 612
rect 1136 614 1138 622
rect 1128 612 1138 614
rect 1136 610 1138 612
rect 1177 614 1179 622
rect 1302 618 1304 624
rect 1392 618 1394 624
rect 1286 616 1289 618
rect 1297 616 1307 618
rect 1376 616 1379 618
rect 1387 616 1397 618
rect 1169 612 1179 614
rect 1177 610 1179 612
rect 136 607 149 609
rect 157 607 160 609
rect 226 607 239 609
rect 247 607 250 609
rect 327 600 329 606
rect 938 608 951 610
rect 959 608 962 610
rect 311 598 314 600
rect 322 598 332 600
rect 116 591 118 597
rect 206 591 208 597
rect 100 589 103 591
rect 111 589 121 591
rect 190 589 193 591
rect 201 589 211 591
rect 326 590 336 592
rect 344 590 347 592
rect 402 594 404 602
rect 852 601 865 603
rect 873 601 876 603
rect 1301 608 1311 610
rect 1319 608 1322 610
rect 1391 608 1401 610
rect 1409 608 1412 610
rect 855 597 857 601
rect 394 592 404 594
rect 402 590 404 592
rect 1018 599 1020 602
rect 1057 599 1059 602
rect 1097 599 1099 602
rect 1136 599 1138 602
rect 1177 599 1179 602
rect 1305 599 1307 608
rect 1395 599 1397 608
rect 918 592 920 598
rect 115 581 125 583
rect 133 581 136 583
rect 205 581 215 583
rect 223 581 226 583
rect 330 581 332 590
rect 795 583 797 591
rect 902 590 905 592
rect 913 590 923 592
rect 119 572 121 581
rect 209 572 211 581
rect 402 579 404 582
rect 782 581 785 583
rect 793 581 805 583
rect 813 581 816 583
rect 917 582 927 584
rect 935 582 938 584
rect 1322 582 1335 584
rect 1343 582 1346 584
rect 1412 582 1425 584
rect 1433 582 1436 584
rect 921 573 923 582
rect 1325 578 1327 582
rect 1006 572 1008 575
rect 1415 578 1417 582
rect 347 564 360 566
rect 368 564 371 566
rect 350 560 352 564
rect 136 555 149 557
rect 157 555 160 557
rect 226 555 239 557
rect 247 555 250 557
rect 855 560 857 564
rect 852 558 865 560
rect 873 558 876 560
rect 139 551 141 555
rect 229 551 231 555
rect 938 556 951 558
rect 959 556 962 558
rect 941 552 943 556
rect 1006 556 1008 564
rect 998 554 1008 556
rect 1006 552 1008 554
rect 832 542 834 548
rect 38 537 40 541
rect 816 540 819 542
rect 827 540 837 542
rect 1006 541 1008 544
rect 35 535 48 537
rect 56 535 59 537
rect 831 532 841 534
rect 849 532 852 534
rect 89 526 91 529
rect 15 519 17 525
rect -1 517 2 519
rect 10 517 20 519
rect 325 521 327 524
rect 835 523 837 532
rect 14 509 24 511
rect 32 509 35 511
rect 18 500 20 509
rect 89 510 91 518
rect 81 508 91 510
rect 89 506 91 508
rect 325 505 327 513
rect 785 509 787 512
rect 1321 510 1323 514
rect 1411 510 1413 514
rect 317 503 327 505
rect 325 501 327 503
rect 1318 508 1331 510
rect 1339 508 1342 510
rect 1408 508 1421 510
rect 1429 508 1432 510
rect 852 506 865 508
rect 873 506 876 508
rect 855 502 857 506
rect 89 495 91 498
rect 325 490 327 493
rect 395 491 397 495
rect 392 489 405 491
rect 413 489 416 491
rect 785 493 787 501
rect 777 491 787 493
rect 1298 492 1300 498
rect 1388 492 1390 498
rect 785 489 787 491
rect 1282 490 1285 492
rect 1293 490 1303 492
rect 1372 490 1375 492
rect 1383 490 1393 492
rect 35 483 48 485
rect 56 483 59 485
rect 38 479 40 483
rect -164 473 -162 476
rect -125 473 -123 476
rect -85 473 -83 476
rect -46 473 -44 476
rect -5 473 -3 476
rect 143 479 145 483
rect 233 479 235 483
rect 1297 482 1307 484
rect 1315 482 1318 484
rect 1387 482 1397 484
rect 1405 482 1408 484
rect 140 477 153 479
rect 161 477 164 479
rect 230 477 243 479
rect 251 477 254 479
rect 372 473 374 479
rect 785 478 787 481
rect 1301 473 1303 482
rect 1391 473 1393 482
rect 356 471 359 473
rect 367 471 377 473
rect -164 457 -162 465
rect -172 455 -162 457
rect -164 453 -162 455
rect -125 457 -123 465
rect -133 455 -123 457
rect -125 453 -123 455
rect -85 457 -83 465
rect -93 455 -83 457
rect -85 453 -83 455
rect -46 457 -44 465
rect -54 455 -44 457
rect -46 453 -44 455
rect -5 457 -3 465
rect 120 461 122 467
rect 210 461 212 467
rect 371 463 381 465
rect 389 463 392 465
rect 104 459 107 461
rect 115 459 125 461
rect 194 459 197 461
rect 205 459 215 461
rect -13 455 -3 457
rect -5 453 -3 455
rect 375 454 377 463
rect 1318 456 1331 458
rect 1339 456 1342 458
rect 1408 456 1421 458
rect 1429 456 1432 458
rect 119 451 129 453
rect 137 451 140 453
rect 209 451 219 453
rect 227 451 230 453
rect -164 442 -162 445
rect -125 442 -123 445
rect -85 442 -83 445
rect -46 442 -44 445
rect -5 442 -3 445
rect 123 442 125 451
rect 213 442 215 451
rect 1321 452 1323 456
rect 481 446 483 450
rect 1411 452 1413 456
rect 478 444 491 446
rect 499 444 502 446
rect 392 437 405 439
rect 413 437 416 439
rect 1220 438 1222 442
rect 395 433 397 437
rect 1217 436 1230 438
rect 1238 436 1241 438
rect 458 428 460 434
rect 140 425 153 427
rect 161 425 164 427
rect 230 425 243 427
rect 251 425 254 427
rect 143 421 145 425
rect -176 415 -174 418
rect 233 421 235 425
rect 335 419 337 427
rect 442 426 445 428
rect 453 426 463 428
rect 1271 427 1273 430
rect 1197 420 1199 426
rect 322 417 325 419
rect 333 417 345 419
rect 353 417 356 419
rect 457 418 467 420
rect 475 418 478 420
rect 1181 418 1184 420
rect 1192 418 1202 420
rect 461 409 463 418
rect 1196 410 1206 412
rect 1214 410 1217 412
rect -176 399 -174 407
rect 1200 401 1202 410
rect 1271 411 1273 419
rect 1263 409 1273 411
rect 1271 407 1273 409
rect -184 397 -174 399
rect -176 395 -174 397
rect 395 396 397 400
rect 392 394 405 396
rect 413 394 416 396
rect 1271 396 1273 399
rect 478 392 491 394
rect 499 392 502 394
rect 481 388 483 392
rect -176 384 -174 387
rect 1217 384 1230 386
rect 1238 384 1241 386
rect 372 378 374 384
rect 1220 380 1222 384
rect 356 376 359 378
rect 367 376 377 378
rect 1018 374 1020 377
rect 1057 374 1059 377
rect 1097 374 1099 377
rect 1136 374 1138 377
rect 1177 374 1179 377
rect 1325 380 1327 384
rect 1415 380 1417 384
rect 1322 378 1335 380
rect 1343 378 1346 380
rect 1412 378 1425 380
rect 1433 378 1436 380
rect 371 368 381 370
rect 389 368 392 370
rect 139 353 141 357
rect 375 359 377 368
rect 229 353 231 357
rect 1018 358 1020 366
rect 1010 356 1020 358
rect 1018 354 1020 356
rect 1057 358 1059 366
rect 1049 356 1059 358
rect 1057 354 1059 356
rect 1097 358 1099 366
rect 1089 356 1099 358
rect 1097 354 1099 356
rect 1136 358 1138 366
rect 1128 356 1138 358
rect 1136 354 1138 356
rect 1177 358 1179 366
rect 1302 362 1304 368
rect 1392 362 1394 368
rect 1286 360 1289 362
rect 1297 360 1307 362
rect 1376 360 1379 362
rect 1387 360 1397 362
rect 1169 356 1179 358
rect 1177 354 1179 356
rect 136 351 149 353
rect 157 351 160 353
rect 226 351 239 353
rect 247 351 250 353
rect 1301 352 1311 354
rect 1319 352 1322 354
rect 1391 352 1401 354
rect 1409 352 1412 354
rect 392 342 405 344
rect 413 342 416 344
rect 1018 343 1020 346
rect 1057 343 1059 346
rect 1097 343 1099 346
rect 1136 343 1138 346
rect 1177 343 1179 346
rect 1305 343 1307 352
rect 1395 343 1397 352
rect 116 335 118 341
rect 206 335 208 341
rect 395 338 397 342
rect 100 333 103 335
rect 111 333 121 335
rect 190 333 193 335
rect 201 333 211 335
rect 115 325 125 327
rect 133 325 136 327
rect 205 325 215 327
rect 223 325 226 327
rect 1322 326 1335 328
rect 1343 326 1346 328
rect 1412 326 1425 328
rect 1433 326 1436 328
rect 119 316 121 325
rect 209 316 211 325
rect 1325 322 1327 326
rect 1006 316 1008 319
rect 1415 322 1417 326
rect 136 299 149 301
rect 157 299 160 301
rect 226 299 239 301
rect 247 299 250 301
rect 139 295 141 299
rect 229 295 231 299
rect 1006 300 1008 308
rect 998 298 1008 300
rect 1006 296 1008 298
rect 38 281 40 285
rect 350 283 352 287
rect 1006 285 1008 288
rect 347 281 360 283
rect 368 281 371 283
rect 35 279 48 281
rect 56 279 59 281
rect 402 275 404 278
rect 89 270 91 273
rect 15 263 17 269
rect -1 261 2 263
rect 10 261 20 263
rect 327 265 329 271
rect 311 263 314 265
rect 322 263 332 265
rect 14 253 24 255
rect 32 253 35 255
rect 18 244 20 253
rect 89 254 91 262
rect 326 255 336 257
rect 344 255 347 257
rect 402 259 404 267
rect 394 257 404 259
rect 402 255 404 257
rect 81 252 91 254
rect 89 250 91 252
rect 330 246 332 255
rect 402 244 404 247
rect 89 239 91 242
rect 35 227 48 229
rect 56 227 59 229
rect 38 223 40 227
rect -164 217 -162 220
rect -125 217 -123 220
rect -85 217 -83 220
rect -46 217 -44 220
rect -5 217 -3 220
rect 143 223 145 227
rect 347 229 360 231
rect 368 229 371 231
rect 233 223 235 227
rect 350 225 352 229
rect 140 221 153 223
rect 161 221 164 223
rect 230 221 243 223
rect 251 221 254 223
rect -164 201 -162 209
rect -172 199 -162 201
rect -164 197 -162 199
rect -125 201 -123 209
rect -133 199 -123 201
rect -125 197 -123 199
rect -85 201 -83 209
rect -93 199 -83 201
rect -85 197 -83 199
rect -46 201 -44 209
rect -54 199 -44 201
rect -46 197 -44 199
rect -5 201 -3 209
rect 120 205 122 211
rect 210 205 212 211
rect 104 203 107 205
rect 115 203 125 205
rect 194 203 197 205
rect 205 203 215 205
rect -13 199 -3 201
rect -5 197 -3 199
rect 119 195 129 197
rect 137 195 140 197
rect 209 195 219 197
rect 227 195 230 197
rect -164 186 -162 189
rect -125 186 -123 189
rect -85 186 -83 189
rect -46 186 -44 189
rect -5 186 -3 189
rect 123 186 125 195
rect 213 186 215 195
rect 140 169 153 171
rect 161 169 164 171
rect 230 169 243 171
rect 251 169 254 171
rect 143 165 145 169
rect -176 159 -174 162
rect 233 165 235 169
rect -176 143 -174 151
rect -184 141 -174 143
rect -176 139 -174 141
rect -176 128 -174 131
rect 139 97 141 101
rect 229 97 231 101
rect 136 95 149 97
rect 157 95 160 97
rect 226 95 239 97
rect 247 95 250 97
rect 116 79 118 85
rect 206 79 208 85
rect 100 77 103 79
rect 111 77 121 79
rect 190 77 193 79
rect 201 77 211 79
rect 115 69 125 71
rect 133 69 136 71
rect 205 69 215 71
rect 223 69 226 71
rect 119 60 121 69
rect 209 60 211 69
rect 136 43 149 45
rect 157 43 160 45
rect 226 43 239 45
rect 247 43 250 45
rect 139 39 141 43
rect 229 39 231 43
rect 38 25 40 29
rect 35 23 48 25
rect 56 23 59 25
rect 89 14 91 17
rect 15 7 17 13
rect -1 5 2 7
rect 10 5 20 7
rect 14 -3 24 -1
rect 32 -3 35 -1
rect 18 -12 20 -3
rect 89 -2 91 6
rect 81 -4 91 -2
rect 89 -6 91 -4
rect 89 -17 91 -14
rect 35 -29 48 -27
rect 56 -29 59 -27
rect 38 -33 40 -29
rect -164 -39 -162 -36
rect -125 -39 -123 -36
rect -85 -39 -83 -36
rect -46 -39 -44 -36
rect -5 -39 -3 -36
rect 143 -33 145 -29
rect 233 -33 235 -29
rect 140 -35 153 -33
rect 161 -35 164 -33
rect 230 -35 243 -33
rect 251 -35 254 -33
rect -164 -55 -162 -47
rect -172 -57 -162 -55
rect -164 -59 -162 -57
rect -125 -55 -123 -47
rect -133 -57 -123 -55
rect -125 -59 -123 -57
rect -85 -55 -83 -47
rect -93 -57 -83 -55
rect -85 -59 -83 -57
rect -46 -55 -44 -47
rect -54 -57 -44 -55
rect -46 -59 -44 -57
rect -5 -55 -3 -47
rect 120 -51 122 -45
rect 210 -51 212 -45
rect 104 -53 107 -51
rect 115 -53 125 -51
rect 194 -53 197 -51
rect 205 -53 215 -51
rect -13 -57 -3 -55
rect -5 -59 -3 -57
rect 119 -61 129 -59
rect 137 -61 140 -59
rect 209 -61 219 -59
rect 227 -61 230 -59
rect -164 -70 -162 -67
rect -125 -70 -123 -67
rect -85 -70 -83 -67
rect -46 -70 -44 -67
rect -5 -70 -3 -67
rect 123 -70 125 -61
rect 213 -70 215 -61
rect 140 -87 153 -85
rect 161 -87 164 -85
rect 230 -87 243 -85
rect 251 -87 254 -85
rect 143 -91 145 -87
rect -176 -97 -174 -94
rect 233 -91 235 -87
rect -176 -113 -174 -105
rect -184 -115 -174 -113
rect -176 -117 -174 -115
rect -176 -128 -174 -125
<< polycontact >>
rect 138 1893 142 1897
rect 228 1893 232 1897
rect 115 1877 119 1881
rect 205 1877 209 1881
rect 118 1848 122 1852
rect 208 1848 212 1852
rect 138 1827 142 1831
rect 228 1827 232 1831
rect 37 1821 41 1825
rect 14 1805 18 1809
rect 77 1787 81 1791
rect 17 1776 21 1780
rect 142 1763 146 1767
rect 37 1755 41 1759
rect 232 1763 236 1767
rect 119 1747 123 1751
rect 209 1747 213 1751
rect -176 1734 -172 1738
rect -137 1734 -133 1738
rect -97 1734 -93 1738
rect -58 1734 -54 1738
rect -17 1734 -13 1738
rect 122 1718 126 1722
rect 212 1718 216 1722
rect 142 1697 146 1701
rect 232 1697 236 1701
rect -188 1676 -184 1680
rect 138 1637 142 1641
rect 228 1637 232 1641
rect 115 1621 119 1625
rect 205 1621 209 1625
rect 118 1592 122 1596
rect 208 1592 212 1596
rect 138 1571 142 1575
rect 228 1571 232 1575
rect 37 1565 41 1569
rect 14 1549 18 1553
rect 77 1531 81 1535
rect 1320 1538 1324 1542
rect 1410 1538 1414 1542
rect 17 1520 21 1524
rect 1297 1522 1301 1526
rect 1387 1522 1391 1526
rect 142 1507 146 1511
rect 37 1499 41 1503
rect 232 1507 236 1511
rect 313 1507 317 1511
rect 394 1500 398 1504
rect 119 1491 123 1495
rect 209 1491 213 1495
rect 1300 1493 1304 1497
rect 1390 1493 1394 1497
rect -176 1478 -172 1482
rect -137 1478 -133 1482
rect -97 1478 -93 1482
rect -58 1478 -54 1482
rect -17 1478 -13 1482
rect 371 1484 375 1488
rect 1320 1472 1324 1476
rect 1410 1472 1414 1476
rect 122 1462 126 1466
rect 212 1462 216 1466
rect 1219 1466 1223 1470
rect 374 1455 378 1459
rect 480 1455 484 1459
rect 1196 1450 1200 1454
rect 142 1441 146 1445
rect 232 1441 236 1445
rect 334 1432 338 1436
rect 394 1434 398 1438
rect 457 1439 461 1443
rect -188 1420 -184 1424
rect 1259 1432 1263 1436
rect 1199 1421 1203 1425
rect 460 1410 464 1414
rect 394 1405 398 1409
rect 1324 1408 1328 1412
rect 1219 1400 1223 1404
rect 1414 1408 1418 1412
rect 371 1389 375 1393
rect 480 1389 484 1393
rect 1301 1392 1305 1396
rect 1391 1392 1395 1396
rect 138 1381 142 1385
rect 228 1381 232 1385
rect 1006 1379 1010 1383
rect 1045 1379 1049 1383
rect 1085 1379 1089 1383
rect 1124 1379 1128 1383
rect 1165 1379 1169 1383
rect 115 1365 119 1369
rect 205 1365 209 1369
rect 773 1365 777 1369
rect 374 1360 378 1364
rect 1304 1363 1308 1367
rect 1394 1363 1398 1367
rect 854 1358 858 1362
rect 118 1336 122 1340
rect 208 1336 212 1340
rect 394 1339 398 1343
rect 831 1342 835 1346
rect 1324 1342 1328 1346
rect 1414 1342 1418 1346
rect 138 1315 142 1319
rect 228 1315 232 1319
rect 994 1321 998 1325
rect 834 1313 838 1317
rect 940 1313 944 1317
rect 37 1309 41 1313
rect 14 1293 18 1297
rect 349 1292 353 1296
rect 794 1290 798 1294
rect 854 1292 858 1296
rect 917 1297 921 1301
rect 77 1275 81 1279
rect 1320 1282 1324 1286
rect 326 1276 330 1280
rect 17 1264 21 1268
rect 1410 1282 1414 1286
rect 390 1261 394 1265
rect 920 1268 924 1272
rect 854 1263 858 1267
rect 1297 1266 1301 1270
rect 1387 1266 1391 1270
rect 142 1251 146 1255
rect 37 1243 41 1247
rect 232 1251 236 1255
rect 329 1247 333 1251
rect 831 1247 835 1251
rect 940 1247 944 1251
rect 119 1235 123 1239
rect 209 1235 213 1239
rect -176 1222 -172 1226
rect -137 1222 -133 1226
rect -97 1222 -93 1226
rect -58 1222 -54 1226
rect -17 1222 -13 1226
rect 1300 1237 1304 1241
rect 1390 1237 1394 1241
rect 349 1226 353 1230
rect 834 1218 838 1222
rect 1320 1216 1324 1220
rect 1410 1216 1414 1220
rect 122 1206 126 1210
rect 212 1206 216 1210
rect 1219 1210 1223 1214
rect 854 1197 858 1201
rect 1196 1194 1200 1198
rect 142 1185 146 1189
rect 232 1185 236 1189
rect -188 1164 -184 1168
rect 313 1172 317 1176
rect 1259 1176 1263 1180
rect 394 1165 398 1169
rect 1199 1165 1203 1169
rect 371 1149 375 1153
rect 1324 1152 1328 1156
rect 138 1125 142 1129
rect 228 1125 232 1129
rect 773 1132 777 1136
rect 1219 1144 1223 1148
rect 1414 1152 1418 1156
rect 1301 1136 1305 1140
rect 1391 1136 1395 1140
rect 374 1120 378 1124
rect 480 1120 484 1124
rect 854 1125 858 1129
rect 1006 1123 1010 1127
rect 1045 1123 1049 1127
rect 1085 1123 1089 1127
rect 1124 1123 1128 1127
rect 1165 1123 1169 1127
rect 115 1109 119 1113
rect 205 1109 209 1113
rect 831 1109 835 1113
rect 334 1097 338 1101
rect 394 1099 398 1103
rect 457 1104 461 1108
rect 1304 1107 1308 1111
rect 1394 1107 1398 1111
rect 118 1080 122 1084
rect 208 1080 212 1084
rect 1324 1086 1328 1090
rect 1414 1086 1418 1090
rect 834 1080 838 1084
rect 940 1080 944 1084
rect 460 1075 464 1079
rect 394 1070 398 1074
rect 138 1059 142 1063
rect 228 1059 232 1063
rect 37 1053 41 1057
rect 371 1054 375 1058
rect 480 1054 484 1058
rect 794 1057 798 1061
rect 854 1059 858 1063
rect 917 1064 921 1068
rect 994 1065 998 1069
rect 14 1037 18 1041
rect 77 1019 81 1023
rect 920 1035 924 1039
rect 374 1025 378 1029
rect 854 1030 858 1034
rect 1320 1026 1324 1030
rect 17 1008 21 1012
rect 539 1012 543 1016
rect 394 1004 398 1008
rect 577 1012 581 1016
rect 615 1012 619 1016
rect 653 1012 657 1016
rect 718 1013 722 1017
rect 1410 1026 1414 1030
rect 831 1014 835 1018
rect 940 1014 944 1018
rect 1297 1010 1301 1014
rect 1387 1010 1391 1014
rect 142 995 146 999
rect 37 987 41 991
rect 232 995 236 999
rect 834 985 838 989
rect 119 979 123 983
rect 209 979 213 983
rect 1300 981 1304 985
rect 1390 981 1394 985
rect -176 966 -172 970
rect -137 966 -133 970
rect -97 966 -93 970
rect -58 966 -54 970
rect -17 966 -13 970
rect 672 976 676 980
rect 702 977 706 981
rect 643 965 647 969
rect 349 957 353 961
rect 122 950 126 954
rect 212 950 216 954
rect 718 956 722 960
rect 854 964 858 968
rect 1320 960 1324 964
rect 1410 960 1414 964
rect 326 941 330 945
rect 142 929 146 933
rect 232 929 236 933
rect 1219 954 1223 958
rect 390 926 394 930
rect 634 935 638 939
rect 1196 938 1200 942
rect -188 908 -184 912
rect 605 924 609 928
rect 329 912 333 916
rect 1259 920 1263 924
rect 349 891 353 895
rect 718 899 722 903
rect 773 899 777 903
rect 1199 909 1203 913
rect 596 894 600 898
rect 1324 896 1328 900
rect 854 892 858 896
rect 567 883 571 887
rect 1219 888 1223 892
rect 1414 896 1418 900
rect 138 869 142 873
rect 228 869 232 873
rect 537 872 541 876
rect 831 876 835 880
rect 1301 880 1305 884
rect 1391 880 1395 884
rect 1006 867 1010 871
rect 1045 867 1049 871
rect 1085 867 1089 871
rect 1124 867 1128 871
rect 1165 867 1169 871
rect 115 853 119 857
rect 205 853 209 857
rect 313 837 317 841
rect 529 843 533 847
rect 718 842 722 846
rect 1304 851 1308 855
rect 1394 851 1398 855
rect 834 847 838 851
rect 940 847 944 851
rect 394 830 398 834
rect 118 824 122 828
rect 208 824 212 828
rect 794 824 798 828
rect 854 826 858 830
rect 917 831 921 835
rect 1324 830 1328 834
rect 1414 830 1418 834
rect 371 814 375 818
rect 521 814 525 818
rect 138 803 142 807
rect 228 803 232 807
rect 994 809 998 813
rect 920 802 924 806
rect 37 797 41 801
rect 854 797 858 801
rect 374 785 378 789
rect 480 785 484 789
rect 14 781 18 785
rect 831 781 835 785
rect 940 781 944 785
rect 77 763 81 767
rect 334 762 338 766
rect 394 764 398 768
rect 457 769 461 773
rect 1320 770 1324 774
rect 1410 770 1414 774
rect 17 752 21 756
rect 834 752 838 756
rect 1297 754 1301 758
rect 1387 754 1391 758
rect 142 739 146 743
rect 37 731 41 735
rect 232 739 236 743
rect 460 740 464 744
rect 394 735 398 739
rect 854 731 858 735
rect 119 723 123 727
rect 209 723 213 727
rect -176 710 -172 714
rect -137 710 -133 714
rect -97 710 -93 714
rect -58 710 -54 714
rect -17 710 -13 714
rect 371 719 375 723
rect 480 719 484 723
rect 1300 725 1304 729
rect 1390 725 1394 729
rect 1320 704 1324 708
rect 1410 704 1414 708
rect 122 694 126 698
rect 212 694 216 698
rect 1219 698 1223 702
rect 374 690 378 694
rect 142 673 146 677
rect 232 673 236 677
rect 1196 682 1200 686
rect 394 669 398 673
rect 773 666 777 670
rect -188 652 -184 656
rect 854 659 858 663
rect 1259 664 1263 668
rect 1199 653 1203 657
rect 831 643 835 647
rect 1324 640 1328 644
rect 1219 632 1223 636
rect 1414 640 1418 644
rect 349 622 353 626
rect 1301 624 1305 628
rect 1391 624 1395 628
rect 138 613 142 617
rect 228 613 232 617
rect 834 614 838 618
rect 940 614 944 618
rect 1006 611 1010 615
rect 1045 611 1049 615
rect 1085 611 1089 615
rect 1124 611 1128 615
rect 1165 611 1169 615
rect 326 606 330 610
rect 115 597 119 601
rect 205 597 209 601
rect 390 591 394 595
rect 794 591 798 595
rect 854 593 858 597
rect 917 598 921 602
rect 1304 595 1308 599
rect 1394 595 1398 599
rect 329 577 333 581
rect 118 568 122 572
rect 208 568 212 572
rect 920 569 924 573
rect 1324 574 1328 578
rect 1414 574 1418 578
rect 854 564 858 568
rect 349 556 353 560
rect 138 547 142 551
rect 228 547 232 551
rect 831 548 835 552
rect 940 548 944 552
rect 994 553 998 557
rect 37 541 41 545
rect 14 525 18 529
rect 77 507 81 511
rect 834 519 838 523
rect 1320 514 1324 518
rect 17 496 21 500
rect 313 502 317 506
rect 1410 514 1414 518
rect 394 495 398 499
rect 773 490 777 494
rect 854 498 858 502
rect 1297 498 1301 502
rect 1387 498 1391 502
rect 142 483 146 487
rect 37 475 41 479
rect 232 483 236 487
rect 371 479 375 483
rect 119 467 123 471
rect 209 467 213 471
rect -176 454 -172 458
rect -137 454 -133 458
rect -97 454 -93 458
rect -58 454 -54 458
rect -17 454 -13 458
rect 1300 469 1304 473
rect 1390 469 1394 473
rect 374 450 378 454
rect 480 450 484 454
rect 1320 448 1324 452
rect 1410 448 1414 452
rect 122 438 126 442
rect 212 438 216 442
rect 1219 442 1223 446
rect 334 427 338 431
rect 394 429 398 433
rect 457 434 461 438
rect 142 417 146 421
rect 232 417 236 421
rect 1196 426 1200 430
rect -188 396 -184 400
rect 460 405 464 409
rect 394 400 398 404
rect 1259 408 1263 412
rect 1199 397 1203 401
rect 371 384 375 388
rect 480 384 484 388
rect 1324 384 1328 388
rect 1219 376 1223 380
rect 1414 384 1418 388
rect 138 357 142 361
rect 228 357 232 361
rect 1301 368 1305 372
rect 1391 368 1395 372
rect 374 355 378 359
rect 1006 355 1010 359
rect 1045 355 1049 359
rect 1085 355 1089 359
rect 1124 355 1128 359
rect 1165 355 1169 359
rect 115 341 119 345
rect 205 341 209 345
rect 394 334 398 338
rect 1304 339 1308 343
rect 1394 339 1398 343
rect 1324 318 1328 322
rect 1414 318 1418 322
rect 118 312 122 316
rect 208 312 212 316
rect 138 291 142 295
rect 228 291 232 295
rect 994 297 998 301
rect 37 285 41 289
rect 349 287 353 291
rect 14 269 18 273
rect 326 271 330 275
rect 77 251 81 255
rect 390 256 394 260
rect 17 240 21 244
rect 329 242 333 246
rect 142 227 146 231
rect 37 219 41 223
rect 232 227 236 231
rect 349 221 353 225
rect 119 211 123 215
rect 209 211 213 215
rect -176 198 -172 202
rect -137 198 -133 202
rect -97 198 -93 202
rect -58 198 -54 202
rect -17 198 -13 202
rect 122 182 126 186
rect 212 182 216 186
rect 142 161 146 165
rect 232 161 236 165
rect -188 140 -184 144
rect 138 101 142 105
rect 228 101 232 105
rect 115 85 119 89
rect 205 85 209 89
rect 118 56 122 60
rect 208 56 212 60
rect 138 35 142 39
rect 228 35 232 39
rect 37 29 41 33
rect 14 13 18 17
rect 77 -5 81 -1
rect 17 -16 21 -12
rect 142 -29 146 -25
rect 37 -37 41 -33
rect 232 -29 236 -25
rect 119 -45 123 -41
rect 209 -45 213 -41
rect -176 -58 -172 -54
rect -137 -58 -133 -54
rect -97 -58 -93 -54
rect -58 -58 -54 -54
rect -17 -58 -13 -54
rect 122 -74 126 -70
rect 212 -74 216 -70
rect 142 -95 146 -91
rect 232 -95 236 -91
rect -188 -116 -184 -112
<< metal1 >>
rect -195 1900 142 1904
rect 174 1900 232 1904
rect -195 1680 -191 1900
rect 115 1881 119 1900
rect 138 1897 142 1900
rect 162 1894 166 1900
rect 157 1890 166 1894
rect 93 1876 97 1880
rect 93 1872 103 1876
rect 93 1860 97 1872
rect 111 1864 125 1868
rect 149 1866 157 1882
rect 162 1875 166 1890
rect 174 1866 178 1900
rect 205 1881 209 1900
rect 228 1897 232 1900
rect 252 1894 256 1900
rect 247 1890 256 1894
rect 149 1862 178 1866
rect 183 1876 187 1880
rect 183 1872 193 1876
rect 149 1860 157 1862
rect 183 1860 187 1872
rect 201 1864 215 1868
rect 239 1866 247 1882
rect 252 1875 256 1890
rect 239 1862 288 1866
rect 239 1860 247 1862
rect 133 1856 157 1860
rect 223 1856 247 1860
rect -183 1833 18 1837
rect -183 1738 -179 1833
rect 14 1832 18 1833
rect 14 1828 41 1832
rect 14 1809 18 1828
rect 37 1825 41 1828
rect 61 1822 65 1828
rect 56 1818 65 1822
rect -8 1804 -4 1808
rect -8 1800 2 1804
rect -8 1788 -4 1800
rect 10 1792 24 1796
rect 48 1791 56 1810
rect 61 1803 65 1818
rect 118 1823 122 1848
rect 149 1842 157 1856
rect 162 1834 166 1849
rect 157 1830 166 1834
rect 138 1823 142 1827
rect 162 1824 166 1830
rect 118 1819 142 1823
rect 208 1823 212 1848
rect 239 1842 247 1856
rect 252 1834 256 1849
rect 247 1830 256 1834
rect 228 1823 232 1827
rect 252 1824 256 1830
rect 208 1819 232 1823
rect 78 1811 102 1815
rect 84 1806 88 1811
rect 92 1791 96 1798
rect 118 1791 122 1819
rect 208 1810 212 1819
rect 208 1806 272 1810
rect 48 1788 77 1791
rect 32 1787 77 1788
rect 92 1787 123 1791
rect 32 1784 56 1787
rect 92 1786 96 1787
rect -175 1758 -151 1762
rect -136 1758 -112 1762
rect -96 1758 -72 1762
rect -57 1758 -33 1762
rect -16 1758 8 1762
rect -169 1753 -165 1758
rect -130 1753 -126 1758
rect -90 1753 -86 1758
rect -51 1753 -47 1758
rect -10 1753 -6 1758
rect -161 1738 -157 1745
rect -122 1738 -118 1745
rect -82 1738 -78 1745
rect -43 1738 -39 1745
rect -2 1738 2 1745
rect 17 1751 21 1776
rect 48 1770 56 1784
rect 61 1762 65 1777
rect 84 1773 88 1778
rect 119 1774 123 1787
rect 80 1769 100 1773
rect 119 1770 146 1774
rect 178 1771 236 1774
rect 56 1758 65 1762
rect 37 1751 41 1755
rect 61 1752 65 1758
rect 17 1747 41 1751
rect 119 1751 123 1770
rect 142 1767 146 1770
rect 166 1764 170 1770
rect 161 1760 170 1764
rect 17 1738 21 1747
rect -183 1734 -176 1738
rect -161 1734 -137 1738
rect -122 1734 -97 1738
rect -82 1734 -58 1738
rect -43 1734 -17 1738
rect -2 1734 21 1738
rect 97 1746 101 1750
rect 97 1742 107 1746
rect -161 1733 -157 1734
rect -122 1733 -118 1734
rect -82 1733 -78 1734
rect -43 1733 -39 1734
rect -2 1733 2 1734
rect 97 1730 101 1742
rect 115 1734 129 1738
rect 153 1735 161 1752
rect 166 1745 170 1760
rect 178 1735 182 1771
rect 209 1770 236 1771
rect 209 1751 213 1770
rect 232 1767 236 1770
rect 256 1764 260 1770
rect 251 1760 260 1764
rect 153 1732 182 1735
rect 187 1746 191 1750
rect 187 1742 197 1746
rect 153 1730 161 1732
rect 187 1730 191 1742
rect 205 1734 219 1738
rect 243 1736 251 1752
rect 256 1745 260 1760
rect 268 1736 272 1806
rect 243 1732 272 1736
rect 243 1730 251 1732
rect 137 1726 161 1730
rect 227 1726 251 1730
rect -169 1720 -165 1725
rect -130 1720 -126 1725
rect -90 1720 -86 1725
rect -51 1720 -47 1725
rect -10 1720 -6 1725
rect -173 1716 -153 1720
rect -134 1716 -114 1720
rect -94 1716 -74 1720
rect -55 1716 -35 1720
rect -14 1716 6 1720
rect -187 1700 -163 1704
rect -181 1695 -177 1700
rect -173 1680 -169 1687
rect 122 1693 126 1718
rect 153 1712 161 1726
rect 166 1704 170 1719
rect 161 1700 170 1704
rect 142 1693 146 1697
rect 166 1694 170 1700
rect 122 1689 146 1693
rect 212 1693 216 1718
rect 243 1712 251 1726
rect 256 1704 260 1719
rect 251 1700 260 1704
rect 232 1693 236 1697
rect 256 1694 260 1700
rect 212 1689 236 1693
rect 122 1680 126 1689
rect -195 1676 -188 1680
rect -173 1676 126 1680
rect 212 1680 216 1689
rect 284 1680 288 1862
rect 212 1676 288 1680
rect -173 1675 -169 1676
rect -181 1662 -177 1667
rect -185 1658 -165 1662
rect -195 1644 142 1648
rect 174 1644 232 1648
rect -195 1424 -191 1644
rect 115 1625 119 1644
rect 138 1641 142 1644
rect 162 1638 166 1644
rect 157 1634 166 1638
rect 93 1620 97 1624
rect 93 1616 103 1620
rect 93 1604 97 1616
rect 111 1608 125 1612
rect 149 1610 157 1626
rect 162 1619 166 1634
rect 174 1610 178 1644
rect 205 1625 209 1644
rect 228 1641 232 1644
rect 252 1638 256 1644
rect 247 1634 256 1638
rect 149 1606 178 1610
rect 183 1620 187 1624
rect 183 1616 193 1620
rect 149 1604 157 1606
rect 183 1604 187 1616
rect 201 1608 215 1612
rect 239 1610 247 1626
rect 252 1619 256 1634
rect 239 1606 288 1610
rect 239 1604 247 1606
rect 133 1600 157 1604
rect 223 1600 247 1604
rect -183 1577 18 1581
rect -183 1482 -179 1577
rect 14 1576 18 1577
rect 14 1572 41 1576
rect 14 1553 18 1572
rect 37 1569 41 1572
rect 61 1566 65 1572
rect 56 1562 65 1566
rect -8 1548 -4 1552
rect -8 1544 2 1548
rect -8 1532 -4 1544
rect 10 1536 24 1540
rect 48 1535 56 1554
rect 61 1547 65 1562
rect 118 1567 122 1592
rect 149 1586 157 1600
rect 162 1578 166 1593
rect 157 1574 166 1578
rect 138 1567 142 1571
rect 162 1568 166 1574
rect 118 1563 142 1567
rect 208 1567 212 1592
rect 239 1586 247 1600
rect 252 1578 256 1593
rect 247 1574 256 1578
rect 228 1567 232 1571
rect 252 1568 256 1574
rect 208 1563 232 1567
rect 78 1555 102 1559
rect 84 1550 88 1555
rect 92 1535 96 1542
rect 118 1535 122 1563
rect 208 1554 212 1563
rect 208 1550 272 1554
rect 48 1532 77 1535
rect 32 1531 77 1532
rect 92 1531 123 1535
rect 32 1528 56 1531
rect 92 1530 96 1531
rect -175 1502 -151 1506
rect -136 1502 -112 1506
rect -96 1502 -72 1506
rect -57 1502 -33 1506
rect -16 1502 8 1506
rect -169 1497 -165 1502
rect -130 1497 -126 1502
rect -90 1497 -86 1502
rect -51 1497 -47 1502
rect -10 1497 -6 1502
rect -161 1482 -157 1489
rect -122 1482 -118 1489
rect -82 1482 -78 1489
rect -43 1482 -39 1489
rect -2 1482 2 1489
rect 17 1495 21 1520
rect 48 1514 56 1528
rect 61 1506 65 1521
rect 84 1517 88 1522
rect 119 1518 123 1531
rect 80 1513 100 1517
rect 119 1514 146 1518
rect 178 1515 236 1518
rect 56 1502 65 1506
rect 37 1495 41 1499
rect 61 1496 65 1502
rect 17 1491 41 1495
rect 119 1495 123 1514
rect 142 1511 146 1514
rect 166 1508 170 1514
rect 161 1504 170 1508
rect 17 1482 21 1491
rect -183 1478 -176 1482
rect -161 1478 -137 1482
rect -122 1478 -97 1482
rect -82 1478 -58 1482
rect -43 1478 -17 1482
rect -2 1478 21 1482
rect 97 1490 101 1494
rect 97 1486 107 1490
rect -161 1477 -157 1478
rect -122 1477 -118 1478
rect -82 1477 -78 1478
rect -43 1477 -39 1478
rect -2 1477 2 1478
rect 97 1474 101 1486
rect 115 1478 129 1482
rect 153 1479 161 1496
rect 166 1489 170 1504
rect 178 1479 182 1515
rect 209 1514 236 1515
rect 209 1495 213 1514
rect 232 1511 236 1514
rect 256 1508 260 1514
rect 251 1504 260 1508
rect 153 1476 182 1479
rect 187 1490 191 1494
rect 187 1486 197 1490
rect 153 1474 161 1476
rect 187 1474 191 1486
rect 205 1478 219 1482
rect 243 1480 251 1496
rect 256 1489 260 1504
rect 268 1480 272 1550
rect 243 1476 272 1480
rect 243 1474 251 1476
rect 137 1470 161 1474
rect 227 1470 251 1474
rect -169 1464 -165 1469
rect -130 1464 -126 1469
rect -90 1464 -86 1469
rect -51 1464 -47 1469
rect -10 1464 -6 1469
rect -173 1460 -153 1464
rect -134 1460 -114 1464
rect -94 1460 -74 1464
rect -55 1460 -35 1464
rect -14 1460 6 1464
rect -187 1444 -163 1448
rect -181 1439 -177 1444
rect -173 1424 -169 1431
rect 122 1437 126 1462
rect 153 1456 161 1470
rect 166 1448 170 1463
rect 161 1444 170 1448
rect 142 1437 146 1441
rect 166 1438 170 1444
rect 122 1433 146 1437
rect 212 1437 216 1462
rect 243 1456 251 1470
rect 256 1448 260 1463
rect 251 1444 260 1448
rect 232 1437 236 1441
rect 256 1438 260 1444
rect 212 1433 236 1437
rect 122 1424 126 1433
rect -195 1420 -188 1424
rect -173 1420 126 1424
rect 212 1424 216 1433
rect 284 1424 288 1606
rect 987 1545 1324 1549
rect 1356 1545 1414 1549
rect 314 1531 338 1535
rect 320 1526 324 1531
rect 328 1511 332 1518
rect 212 1420 288 1424
rect 304 1507 313 1511
rect 328 1507 398 1511
rect -173 1419 -169 1420
rect -181 1406 -177 1411
rect -185 1402 -165 1406
rect -195 1388 142 1392
rect 174 1388 232 1392
rect -195 1168 -191 1388
rect 115 1369 119 1388
rect 138 1385 142 1388
rect 162 1382 166 1388
rect 157 1378 166 1382
rect 93 1364 97 1368
rect 93 1360 103 1364
rect 93 1348 97 1360
rect 111 1352 125 1356
rect 149 1354 157 1370
rect 162 1363 166 1378
rect 174 1354 178 1388
rect 205 1369 209 1388
rect 228 1385 232 1388
rect 252 1382 256 1388
rect 247 1378 256 1382
rect 149 1350 178 1354
rect 183 1364 187 1368
rect 183 1360 193 1364
rect 149 1348 157 1350
rect 183 1348 187 1360
rect 201 1352 215 1356
rect 239 1354 247 1370
rect 252 1363 256 1378
rect 239 1350 288 1354
rect 239 1348 247 1350
rect 133 1344 157 1348
rect 223 1344 247 1348
rect -183 1321 18 1325
rect -183 1226 -179 1321
rect 14 1320 18 1321
rect 14 1316 41 1320
rect 14 1297 18 1316
rect 37 1313 41 1316
rect 61 1310 65 1316
rect 56 1306 65 1310
rect -8 1292 -4 1296
rect -8 1288 2 1292
rect -8 1276 -4 1288
rect 10 1280 24 1284
rect 48 1279 56 1298
rect 61 1291 65 1306
rect 118 1311 122 1336
rect 149 1330 157 1344
rect 162 1322 166 1337
rect 157 1318 166 1322
rect 138 1311 142 1315
rect 162 1312 166 1318
rect 118 1307 142 1311
rect 208 1311 212 1336
rect 239 1330 247 1344
rect 252 1322 256 1337
rect 247 1318 256 1322
rect 228 1311 232 1315
rect 252 1312 256 1318
rect 208 1307 232 1311
rect 78 1299 102 1303
rect 84 1294 88 1299
rect 92 1279 96 1286
rect 118 1279 122 1307
rect 208 1298 212 1307
rect 208 1294 272 1298
rect 48 1276 77 1279
rect 32 1275 77 1276
rect 92 1275 123 1279
rect 32 1272 56 1275
rect 92 1274 96 1275
rect -175 1246 -151 1250
rect -136 1246 -112 1250
rect -96 1246 -72 1250
rect -57 1246 -33 1250
rect -16 1246 8 1250
rect -169 1241 -165 1246
rect -130 1241 -126 1246
rect -90 1241 -86 1246
rect -51 1241 -47 1246
rect -10 1241 -6 1246
rect -161 1226 -157 1233
rect -122 1226 -118 1233
rect -82 1226 -78 1233
rect -43 1226 -39 1233
rect -2 1226 2 1233
rect 17 1239 21 1264
rect 48 1258 56 1272
rect 61 1250 65 1265
rect 84 1261 88 1266
rect 119 1262 123 1275
rect 80 1257 100 1261
rect 119 1258 146 1262
rect 178 1259 236 1262
rect 56 1246 65 1250
rect 37 1239 41 1243
rect 61 1240 65 1246
rect 17 1235 41 1239
rect 119 1239 123 1258
rect 142 1255 146 1258
rect 166 1252 170 1258
rect 161 1248 170 1252
rect 17 1226 21 1235
rect -183 1222 -176 1226
rect -161 1222 -137 1226
rect -122 1222 -97 1226
rect -82 1222 -58 1226
rect -43 1222 -17 1226
rect -2 1222 21 1226
rect 97 1234 101 1238
rect 97 1230 107 1234
rect -161 1221 -157 1222
rect -122 1221 -118 1222
rect -82 1221 -78 1222
rect -43 1221 -39 1222
rect -2 1221 2 1222
rect 97 1218 101 1230
rect 115 1222 129 1226
rect 153 1223 161 1240
rect 166 1233 170 1248
rect 178 1223 182 1259
rect 209 1258 236 1259
rect 209 1239 213 1258
rect 232 1255 236 1258
rect 256 1252 260 1258
rect 251 1248 260 1252
rect 153 1220 182 1223
rect 187 1234 191 1238
rect 187 1230 197 1234
rect 153 1218 161 1220
rect 187 1218 191 1230
rect 205 1222 219 1226
rect 243 1224 251 1240
rect 256 1233 260 1248
rect 268 1224 272 1294
rect 243 1220 272 1224
rect 243 1218 251 1220
rect 137 1214 161 1218
rect 227 1214 251 1218
rect -169 1208 -165 1213
rect -130 1208 -126 1213
rect -90 1208 -86 1213
rect -51 1208 -47 1213
rect -10 1208 -6 1213
rect -173 1204 -153 1208
rect -134 1204 -114 1208
rect -94 1204 -74 1208
rect -55 1204 -35 1208
rect -14 1204 6 1208
rect -187 1188 -163 1192
rect -181 1183 -177 1188
rect -173 1168 -169 1175
rect 122 1181 126 1206
rect 153 1200 161 1214
rect 166 1192 170 1207
rect 161 1188 170 1192
rect 142 1181 146 1185
rect 166 1182 170 1188
rect 122 1177 146 1181
rect 212 1181 216 1206
rect 243 1200 251 1214
rect 256 1192 260 1207
rect 251 1188 260 1192
rect 232 1181 236 1185
rect 256 1182 260 1188
rect 212 1177 236 1181
rect 122 1168 126 1177
rect -195 1164 -188 1168
rect -173 1164 126 1168
rect 212 1168 216 1177
rect 284 1168 288 1350
rect 304 1335 308 1507
rect 328 1506 332 1507
rect 320 1493 324 1498
rect 316 1489 336 1493
rect 371 1488 375 1507
rect 394 1504 398 1507
rect 418 1501 422 1507
rect 413 1497 422 1501
rect 349 1483 353 1487
rect 349 1479 359 1483
rect 349 1467 353 1479
rect 367 1471 381 1475
rect 405 1473 413 1489
rect 418 1482 422 1497
rect 405 1469 461 1473
rect 405 1467 413 1469
rect 389 1463 413 1467
rect 374 1444 378 1455
rect 405 1449 413 1463
rect 457 1466 461 1469
rect 457 1462 484 1466
rect 334 1440 378 1444
rect 418 1441 422 1456
rect 457 1443 461 1462
rect 480 1459 484 1462
rect 504 1456 508 1462
rect 499 1452 508 1456
rect 334 1436 338 1440
rect 316 1429 320 1433
rect 358 1429 362 1435
rect 316 1425 325 1429
rect 353 1425 362 1429
rect 374 1430 378 1440
rect 413 1437 422 1441
rect 394 1430 398 1434
rect 418 1431 422 1437
rect 435 1438 439 1442
rect 435 1434 445 1438
rect 374 1426 398 1430
rect 316 1413 320 1425
rect 333 1417 345 1421
rect 334 1406 338 1417
rect 358 1411 362 1425
rect 435 1422 439 1434
rect 453 1426 467 1430
rect 491 1428 499 1444
rect 504 1437 508 1452
rect 491 1424 514 1428
rect 491 1422 499 1424
rect 475 1418 499 1422
rect 371 1412 398 1416
rect 371 1406 375 1412
rect 334 1402 375 1406
rect 394 1409 398 1412
rect 418 1406 422 1412
rect 413 1402 422 1406
rect 371 1393 375 1402
rect 349 1388 353 1392
rect 349 1384 359 1388
rect 349 1372 353 1384
rect 367 1376 381 1380
rect 405 1378 413 1394
rect 418 1387 422 1402
rect 460 1385 464 1410
rect 491 1404 499 1418
rect 504 1396 508 1411
rect 499 1392 508 1396
rect 480 1385 484 1389
rect 504 1386 508 1392
rect 774 1389 798 1393
rect 460 1381 484 1385
rect 780 1384 784 1389
rect 460 1378 464 1381
rect 405 1374 464 1378
rect 405 1372 413 1374
rect 389 1368 413 1372
rect 788 1369 792 1376
rect 374 1335 378 1360
rect 405 1354 413 1368
rect 764 1365 773 1369
rect 788 1365 858 1369
rect 418 1346 422 1361
rect 413 1342 422 1346
rect 394 1335 398 1339
rect 418 1336 422 1342
rect 304 1331 398 1335
rect 326 1299 353 1303
rect 326 1280 330 1299
rect 349 1296 353 1299
rect 373 1293 377 1299
rect 368 1289 377 1293
rect 304 1275 308 1279
rect 304 1271 314 1275
rect 304 1259 308 1271
rect 322 1263 336 1267
rect 360 1265 368 1281
rect 373 1274 377 1289
rect 391 1285 415 1289
rect 397 1280 401 1285
rect 405 1265 409 1272
rect 360 1261 390 1265
rect 405 1261 426 1265
rect 360 1259 368 1261
rect 405 1260 409 1261
rect 344 1255 368 1259
rect 329 1222 333 1247
rect 360 1241 368 1255
rect 373 1233 377 1248
rect 397 1247 401 1252
rect 393 1243 413 1247
rect 368 1229 377 1233
rect 349 1222 353 1226
rect 373 1223 377 1229
rect 329 1218 353 1222
rect 314 1196 338 1200
rect 320 1191 324 1196
rect 764 1193 768 1365
rect 788 1364 792 1365
rect 780 1351 784 1356
rect 776 1347 796 1351
rect 831 1346 835 1365
rect 854 1362 858 1365
rect 878 1359 882 1365
rect 873 1355 882 1359
rect 809 1341 813 1345
rect 809 1337 819 1341
rect 809 1325 813 1337
rect 827 1329 841 1333
rect 865 1331 873 1347
rect 878 1340 882 1355
rect 865 1327 921 1331
rect 865 1325 873 1327
rect 849 1321 873 1325
rect 834 1302 838 1313
rect 865 1307 873 1321
rect 917 1324 921 1327
rect 987 1325 991 1545
rect 1297 1526 1301 1545
rect 1320 1542 1324 1545
rect 1344 1539 1348 1545
rect 1339 1535 1348 1539
rect 1275 1521 1279 1525
rect 1275 1517 1285 1521
rect 1275 1505 1279 1517
rect 1293 1509 1307 1513
rect 1331 1511 1339 1527
rect 1344 1520 1348 1535
rect 1356 1511 1360 1545
rect 1387 1526 1391 1545
rect 1410 1542 1414 1545
rect 1434 1539 1438 1545
rect 1429 1535 1438 1539
rect 1331 1507 1360 1511
rect 1365 1521 1369 1525
rect 1365 1517 1375 1521
rect 1331 1505 1339 1507
rect 1365 1505 1369 1517
rect 1383 1509 1397 1513
rect 1421 1511 1429 1527
rect 1434 1520 1438 1535
rect 1421 1507 1470 1511
rect 1421 1505 1429 1507
rect 1315 1501 1339 1505
rect 1405 1501 1429 1505
rect 999 1478 1200 1482
rect 999 1383 1003 1478
rect 1196 1477 1200 1478
rect 1196 1473 1223 1477
rect 1196 1454 1200 1473
rect 1219 1470 1223 1473
rect 1243 1467 1247 1473
rect 1238 1463 1247 1467
rect 1174 1449 1178 1453
rect 1174 1445 1184 1449
rect 1174 1433 1178 1445
rect 1192 1437 1206 1441
rect 1230 1436 1238 1455
rect 1243 1448 1247 1463
rect 1300 1468 1304 1493
rect 1331 1487 1339 1501
rect 1344 1479 1348 1494
rect 1339 1475 1348 1479
rect 1320 1468 1324 1472
rect 1344 1469 1348 1475
rect 1300 1464 1324 1468
rect 1390 1468 1394 1493
rect 1421 1487 1429 1501
rect 1434 1479 1438 1494
rect 1429 1475 1438 1479
rect 1410 1468 1414 1472
rect 1434 1469 1438 1475
rect 1390 1464 1414 1468
rect 1260 1456 1284 1460
rect 1266 1451 1270 1456
rect 1274 1436 1278 1443
rect 1300 1436 1304 1464
rect 1390 1455 1394 1464
rect 1390 1451 1454 1455
rect 1230 1433 1259 1436
rect 1214 1432 1259 1433
rect 1274 1432 1305 1436
rect 1214 1429 1238 1432
rect 1274 1431 1278 1432
rect 1007 1403 1031 1407
rect 1046 1403 1070 1407
rect 1086 1403 1110 1407
rect 1125 1403 1149 1407
rect 1166 1403 1190 1407
rect 1013 1398 1017 1403
rect 1052 1398 1056 1403
rect 1092 1398 1096 1403
rect 1131 1398 1135 1403
rect 1172 1398 1176 1403
rect 1021 1383 1025 1390
rect 1060 1383 1064 1390
rect 1100 1383 1104 1390
rect 1139 1383 1143 1390
rect 1180 1383 1184 1390
rect 1199 1396 1203 1421
rect 1230 1415 1238 1429
rect 1243 1407 1247 1422
rect 1266 1418 1270 1423
rect 1301 1419 1305 1432
rect 1262 1414 1282 1418
rect 1301 1415 1328 1419
rect 1360 1416 1418 1419
rect 1238 1403 1247 1407
rect 1219 1396 1223 1400
rect 1243 1397 1247 1403
rect 1199 1392 1223 1396
rect 1301 1396 1305 1415
rect 1324 1412 1328 1415
rect 1348 1409 1352 1415
rect 1343 1405 1352 1409
rect 1199 1383 1203 1392
rect 999 1379 1006 1383
rect 1021 1379 1045 1383
rect 1060 1379 1085 1383
rect 1100 1379 1124 1383
rect 1139 1379 1165 1383
rect 1180 1379 1203 1383
rect 1279 1391 1283 1395
rect 1279 1387 1289 1391
rect 1021 1378 1025 1379
rect 1060 1378 1064 1379
rect 1100 1378 1104 1379
rect 1139 1378 1143 1379
rect 1180 1378 1184 1379
rect 1279 1375 1283 1387
rect 1297 1379 1311 1383
rect 1335 1380 1343 1397
rect 1348 1390 1352 1405
rect 1360 1380 1364 1416
rect 1391 1415 1418 1416
rect 1391 1396 1395 1415
rect 1414 1412 1418 1415
rect 1438 1409 1442 1415
rect 1433 1405 1442 1409
rect 1335 1377 1364 1380
rect 1369 1391 1373 1395
rect 1369 1387 1379 1391
rect 1335 1375 1343 1377
rect 1369 1375 1373 1387
rect 1387 1379 1401 1383
rect 1425 1381 1433 1397
rect 1438 1390 1442 1405
rect 1450 1381 1454 1451
rect 1425 1377 1454 1381
rect 1425 1375 1433 1377
rect 1319 1371 1343 1375
rect 1409 1371 1433 1375
rect 1013 1365 1017 1370
rect 1052 1365 1056 1370
rect 1092 1365 1096 1370
rect 1131 1365 1135 1370
rect 1172 1365 1176 1370
rect 1009 1361 1029 1365
rect 1048 1361 1068 1365
rect 1088 1361 1108 1365
rect 1127 1361 1147 1365
rect 1168 1361 1188 1365
rect 995 1345 1019 1349
rect 1001 1340 1005 1345
rect 1009 1325 1013 1332
rect 1304 1338 1308 1363
rect 1335 1357 1343 1371
rect 1348 1349 1352 1364
rect 1343 1345 1352 1349
rect 1324 1338 1328 1342
rect 1348 1339 1352 1345
rect 1304 1334 1328 1338
rect 1394 1338 1398 1363
rect 1425 1357 1433 1371
rect 1438 1349 1442 1364
rect 1433 1345 1442 1349
rect 1414 1338 1418 1342
rect 1438 1339 1442 1345
rect 1394 1334 1418 1338
rect 1304 1325 1308 1334
rect 917 1320 944 1324
rect 987 1321 994 1325
rect 1009 1321 1308 1325
rect 1394 1325 1398 1334
rect 1466 1325 1470 1507
rect 1394 1321 1470 1325
rect 1009 1320 1013 1321
rect 794 1298 838 1302
rect 878 1299 882 1314
rect 917 1301 921 1320
rect 940 1317 944 1320
rect 964 1314 968 1320
rect 959 1310 968 1314
rect 794 1294 798 1298
rect 776 1287 780 1291
rect 818 1287 822 1293
rect 776 1283 785 1287
rect 813 1283 822 1287
rect 834 1288 838 1298
rect 873 1295 882 1299
rect 854 1288 858 1292
rect 878 1289 882 1295
rect 895 1296 899 1300
rect 895 1292 905 1296
rect 834 1284 858 1288
rect 776 1271 780 1283
rect 793 1275 805 1279
rect 794 1264 798 1275
rect 818 1269 822 1283
rect 895 1280 899 1292
rect 913 1284 927 1288
rect 951 1286 959 1302
rect 964 1295 968 1310
rect 1001 1307 1005 1312
rect 997 1303 1017 1307
rect 987 1289 1324 1293
rect 1356 1289 1414 1293
rect 951 1282 971 1286
rect 951 1280 959 1282
rect 935 1276 959 1280
rect 831 1270 858 1274
rect 831 1264 835 1270
rect 794 1260 835 1264
rect 854 1267 858 1270
rect 878 1264 882 1270
rect 873 1260 882 1264
rect 831 1251 835 1260
rect 809 1246 813 1250
rect 809 1242 819 1246
rect 809 1230 813 1242
rect 827 1234 841 1238
rect 865 1236 873 1252
rect 878 1245 882 1260
rect 920 1243 924 1268
rect 951 1262 959 1276
rect 964 1254 968 1269
rect 959 1250 968 1254
rect 940 1243 944 1247
rect 964 1244 968 1250
rect 920 1239 944 1243
rect 920 1236 924 1239
rect 865 1232 924 1236
rect 865 1230 873 1232
rect 849 1226 873 1230
rect 834 1193 838 1218
rect 865 1212 873 1226
rect 878 1204 882 1219
rect 873 1200 882 1204
rect 854 1193 858 1197
rect 878 1194 882 1200
rect 764 1189 858 1193
rect 328 1176 332 1183
rect 212 1164 288 1168
rect 304 1172 313 1176
rect 328 1172 398 1176
rect -173 1163 -169 1164
rect -181 1150 -177 1155
rect -185 1146 -165 1150
rect -195 1132 142 1136
rect 174 1132 232 1136
rect -195 912 -191 1132
rect 115 1113 119 1132
rect 138 1129 142 1132
rect 162 1126 166 1132
rect 157 1122 166 1126
rect 93 1108 97 1112
rect 93 1104 103 1108
rect 93 1092 97 1104
rect 111 1096 125 1100
rect 149 1098 157 1114
rect 162 1107 166 1122
rect 174 1098 178 1132
rect 205 1113 209 1132
rect 228 1129 232 1132
rect 252 1126 256 1132
rect 247 1122 256 1126
rect 149 1094 178 1098
rect 183 1108 187 1112
rect 183 1104 193 1108
rect 149 1092 157 1094
rect 183 1092 187 1104
rect 201 1096 215 1100
rect 239 1098 247 1114
rect 252 1107 256 1122
rect 239 1094 288 1098
rect 239 1092 247 1094
rect 133 1088 157 1092
rect 223 1088 247 1092
rect -183 1065 18 1069
rect -183 970 -179 1065
rect 14 1064 18 1065
rect 14 1060 41 1064
rect 14 1041 18 1060
rect 37 1057 41 1060
rect 61 1054 65 1060
rect 56 1050 65 1054
rect -8 1036 -4 1040
rect -8 1032 2 1036
rect -8 1020 -4 1032
rect 10 1024 24 1028
rect 48 1023 56 1042
rect 61 1035 65 1050
rect 118 1055 122 1080
rect 149 1074 157 1088
rect 162 1066 166 1081
rect 157 1062 166 1066
rect 138 1055 142 1059
rect 162 1056 166 1062
rect 118 1051 142 1055
rect 208 1055 212 1080
rect 239 1074 247 1088
rect 252 1066 256 1081
rect 247 1062 256 1066
rect 228 1055 232 1059
rect 252 1056 256 1062
rect 208 1051 232 1055
rect 78 1043 102 1047
rect 84 1038 88 1043
rect 92 1023 96 1030
rect 118 1023 122 1051
rect 208 1042 212 1051
rect 208 1038 272 1042
rect 48 1020 77 1023
rect 32 1019 77 1020
rect 92 1019 123 1023
rect 32 1016 56 1019
rect 92 1018 96 1019
rect -175 990 -151 994
rect -136 990 -112 994
rect -96 990 -72 994
rect -57 990 -33 994
rect -16 990 8 994
rect -169 985 -165 990
rect -130 985 -126 990
rect -90 985 -86 990
rect -51 985 -47 990
rect -10 985 -6 990
rect -161 970 -157 977
rect -122 970 -118 977
rect -82 970 -78 977
rect -43 970 -39 977
rect -2 970 2 977
rect 17 983 21 1008
rect 48 1002 56 1016
rect 61 994 65 1009
rect 84 1005 88 1010
rect 119 1006 123 1019
rect 80 1001 100 1005
rect 119 1002 146 1006
rect 178 1003 236 1006
rect 56 990 65 994
rect 37 983 41 987
rect 61 984 65 990
rect 17 979 41 983
rect 119 983 123 1002
rect 142 999 146 1002
rect 166 996 170 1002
rect 161 992 170 996
rect 17 970 21 979
rect -183 966 -176 970
rect -161 966 -137 970
rect -122 966 -97 970
rect -82 966 -58 970
rect -43 966 -17 970
rect -2 966 21 970
rect 97 978 101 982
rect 97 974 107 978
rect -161 965 -157 966
rect -122 965 -118 966
rect -82 965 -78 966
rect -43 965 -39 966
rect -2 965 2 966
rect 97 962 101 974
rect 115 966 129 970
rect 153 967 161 984
rect 166 977 170 992
rect 178 967 182 1003
rect 209 1002 236 1003
rect 209 983 213 1002
rect 232 999 236 1002
rect 256 996 260 1002
rect 251 992 260 996
rect 153 964 182 967
rect 187 978 191 982
rect 187 974 197 978
rect 153 962 161 964
rect 187 962 191 974
rect 205 966 219 970
rect 243 968 251 984
rect 256 977 260 992
rect 268 968 272 1038
rect 243 964 272 968
rect 243 962 251 964
rect 137 958 161 962
rect 227 958 251 962
rect -169 952 -165 957
rect -130 952 -126 957
rect -90 952 -86 957
rect -51 952 -47 957
rect -10 952 -6 957
rect -173 948 -153 952
rect -134 948 -114 952
rect -94 948 -74 952
rect -55 948 -35 952
rect -14 948 6 952
rect -187 932 -163 936
rect -181 927 -177 932
rect -173 912 -169 919
rect 122 925 126 950
rect 153 944 161 958
rect 166 936 170 951
rect 161 932 170 936
rect 142 925 146 929
rect 166 926 170 932
rect 122 921 146 925
rect 212 925 216 950
rect 243 944 251 958
rect 256 936 260 951
rect 251 932 260 936
rect 232 925 236 929
rect 256 926 260 932
rect 212 921 236 925
rect 122 912 126 921
rect -195 908 -188 912
rect -173 908 126 912
rect 212 912 216 921
rect 284 912 288 1094
rect 304 1000 308 1172
rect 328 1171 332 1172
rect 320 1158 324 1163
rect 316 1154 336 1158
rect 371 1153 375 1172
rect 394 1169 398 1172
rect 418 1166 422 1172
rect 413 1162 422 1166
rect 349 1148 353 1152
rect 349 1144 359 1148
rect 349 1132 353 1144
rect 367 1136 381 1140
rect 405 1138 413 1154
rect 418 1147 422 1162
rect 774 1156 798 1160
rect 780 1151 784 1156
rect 405 1134 461 1138
rect 788 1136 792 1143
rect 405 1132 413 1134
rect 389 1128 413 1132
rect 374 1109 378 1120
rect 405 1114 413 1128
rect 457 1131 461 1134
rect 764 1132 773 1136
rect 788 1132 858 1136
rect 457 1127 484 1131
rect 334 1105 378 1109
rect 418 1106 422 1121
rect 457 1108 461 1127
rect 480 1124 484 1127
rect 504 1121 508 1127
rect 499 1117 508 1121
rect 334 1101 338 1105
rect 316 1094 320 1098
rect 358 1094 362 1100
rect 316 1090 325 1094
rect 353 1090 362 1094
rect 374 1095 378 1105
rect 413 1102 422 1106
rect 394 1095 398 1099
rect 418 1096 422 1102
rect 435 1103 439 1107
rect 435 1099 445 1103
rect 374 1091 398 1095
rect 316 1078 320 1090
rect 333 1082 345 1086
rect 334 1071 338 1082
rect 358 1076 362 1090
rect 435 1087 439 1099
rect 453 1091 467 1095
rect 491 1093 499 1109
rect 504 1102 508 1117
rect 491 1089 514 1093
rect 491 1087 499 1089
rect 475 1083 499 1087
rect 371 1077 398 1081
rect 371 1071 375 1077
rect 334 1067 375 1071
rect 394 1074 398 1077
rect 418 1071 422 1077
rect 413 1067 422 1071
rect 371 1058 375 1067
rect 349 1053 353 1057
rect 349 1049 359 1053
rect 349 1037 353 1049
rect 367 1041 381 1045
rect 405 1043 413 1059
rect 418 1052 422 1067
rect 460 1050 464 1075
rect 491 1069 499 1083
rect 504 1061 508 1076
rect 499 1057 508 1061
rect 480 1050 484 1054
rect 504 1051 508 1057
rect 460 1046 484 1050
rect 527 1047 645 1051
rect 460 1043 464 1046
rect 405 1039 464 1043
rect 405 1037 413 1039
rect 389 1033 413 1037
rect 374 1000 378 1025
rect 405 1019 413 1033
rect 418 1011 422 1026
rect 527 1016 531 1047
rect 536 1036 560 1040
rect 542 1031 546 1036
rect 413 1007 422 1011
rect 394 1000 398 1004
rect 418 1001 422 1007
rect 513 1012 539 1016
rect 304 996 398 1000
rect 326 964 353 968
rect 326 945 330 964
rect 349 961 353 964
rect 373 958 377 964
rect 368 954 377 958
rect 304 940 308 944
rect 304 936 314 940
rect 304 924 308 936
rect 322 928 336 932
rect 360 930 368 946
rect 373 939 377 954
rect 391 950 415 954
rect 397 945 401 950
rect 405 930 409 937
rect 360 926 390 930
rect 405 926 426 930
rect 360 924 368 926
rect 405 925 409 926
rect 344 920 368 924
rect 212 908 288 912
rect -173 907 -169 908
rect -181 894 -177 899
rect -185 890 -165 894
rect 329 887 333 912
rect 360 906 368 920
rect 373 898 377 913
rect 397 912 401 917
rect 393 908 413 912
rect 368 894 377 898
rect 349 887 353 891
rect 373 888 377 894
rect 329 883 353 887
rect -195 876 142 880
rect 174 876 232 880
rect -195 656 -191 876
rect 115 857 119 876
rect 138 873 142 876
rect 162 870 166 876
rect 157 866 166 870
rect 93 852 97 856
rect 93 848 103 852
rect 93 836 97 848
rect 111 840 125 844
rect 149 842 157 858
rect 162 851 166 866
rect 174 842 178 876
rect 205 857 209 876
rect 228 873 232 876
rect 252 870 256 876
rect 247 866 256 870
rect 149 838 178 842
rect 183 852 187 856
rect 183 848 193 852
rect 149 836 157 838
rect 183 836 187 848
rect 201 840 215 844
rect 239 842 247 858
rect 252 851 256 866
rect 314 861 338 865
rect 320 856 324 861
rect 239 838 288 842
rect 328 841 332 848
rect 239 836 247 838
rect 133 832 157 836
rect 223 832 247 836
rect -183 809 18 813
rect -183 714 -179 809
rect 14 808 18 809
rect 14 804 41 808
rect 14 785 18 804
rect 37 801 41 804
rect 61 798 65 804
rect 56 794 65 798
rect -8 780 -4 784
rect -8 776 2 780
rect -8 764 -4 776
rect 10 768 24 772
rect 48 767 56 786
rect 61 779 65 794
rect 118 799 122 824
rect 149 818 157 832
rect 162 810 166 825
rect 157 806 166 810
rect 138 799 142 803
rect 162 800 166 806
rect 118 795 142 799
rect 208 799 212 824
rect 239 818 247 832
rect 252 810 256 825
rect 247 806 256 810
rect 228 799 232 803
rect 252 800 256 806
rect 208 795 232 799
rect 78 787 102 791
rect 84 782 88 787
rect 92 767 96 774
rect 118 767 122 795
rect 208 786 212 795
rect 208 782 272 786
rect 48 764 77 767
rect 32 763 77 764
rect 92 763 123 767
rect 32 760 56 763
rect 92 762 96 763
rect -175 734 -151 738
rect -136 734 -112 738
rect -96 734 -72 738
rect -57 734 -33 738
rect -16 734 8 738
rect -169 729 -165 734
rect -130 729 -126 734
rect -90 729 -86 734
rect -51 729 -47 734
rect -10 729 -6 734
rect -161 714 -157 721
rect -122 714 -118 721
rect -82 714 -78 721
rect -43 714 -39 721
rect -2 714 2 721
rect 17 727 21 752
rect 48 746 56 760
rect 61 738 65 753
rect 84 749 88 754
rect 119 750 123 763
rect 80 745 100 749
rect 119 746 146 750
rect 178 747 236 750
rect 56 734 65 738
rect 37 727 41 731
rect 61 728 65 734
rect 17 723 41 727
rect 119 727 123 746
rect 142 743 146 746
rect 166 740 170 746
rect 161 736 170 740
rect 17 714 21 723
rect -183 710 -176 714
rect -161 710 -137 714
rect -122 710 -97 714
rect -82 710 -58 714
rect -43 710 -17 714
rect -2 710 21 714
rect 97 722 101 726
rect 97 718 107 722
rect -161 709 -157 710
rect -122 709 -118 710
rect -82 709 -78 710
rect -43 709 -39 710
rect -2 709 2 710
rect 97 706 101 718
rect 115 710 129 714
rect 153 711 161 728
rect 166 721 170 736
rect 178 711 182 747
rect 209 746 236 747
rect 209 727 213 746
rect 232 743 236 746
rect 256 740 260 746
rect 251 736 260 740
rect 153 708 182 711
rect 187 722 191 726
rect 187 718 197 722
rect 153 706 161 708
rect 187 706 191 718
rect 205 710 219 714
rect 243 712 251 728
rect 256 721 260 736
rect 268 712 272 782
rect 243 708 272 712
rect 243 706 251 708
rect 137 702 161 706
rect 227 702 251 706
rect -169 696 -165 701
rect -130 696 -126 701
rect -90 696 -86 701
rect -51 696 -47 701
rect -10 696 -6 701
rect -173 692 -153 696
rect -134 692 -114 696
rect -94 692 -74 696
rect -55 692 -35 696
rect -14 692 6 696
rect -187 676 -163 680
rect -181 671 -177 676
rect -173 656 -169 663
rect 122 669 126 694
rect 153 688 161 702
rect 166 680 170 695
rect 161 676 170 680
rect 142 669 146 673
rect 166 670 170 676
rect 122 665 146 669
rect 212 669 216 694
rect 243 688 251 702
rect 256 680 260 695
rect 251 676 260 680
rect 232 669 236 673
rect 256 670 260 676
rect 212 665 236 669
rect 122 656 126 665
rect -195 652 -188 656
rect -173 652 126 656
rect 212 656 216 665
rect 284 656 288 838
rect 304 837 313 841
rect 328 837 398 841
rect 304 665 308 837
rect 328 836 332 837
rect 320 823 324 828
rect 316 819 336 823
rect 371 818 375 837
rect 394 834 398 837
rect 418 831 422 837
rect 413 827 422 831
rect 349 813 353 817
rect 349 809 359 813
rect 349 797 353 809
rect 367 801 381 805
rect 405 803 413 819
rect 418 812 422 827
rect 513 818 517 1012
rect 550 897 554 1023
rect 565 1016 569 1047
rect 574 1036 598 1040
rect 580 1031 584 1036
rect 565 1012 577 1016
rect 588 938 592 1023
rect 603 1016 607 1047
rect 612 1036 636 1040
rect 618 1031 622 1036
rect 603 1012 615 1016
rect 626 979 630 1023
rect 641 1016 645 1047
rect 650 1036 674 1040
rect 719 1037 743 1041
rect 656 1031 660 1036
rect 725 1032 729 1037
rect 641 1012 653 1016
rect 664 1004 668 1023
rect 733 1017 737 1024
rect 712 1013 718 1017
rect 733 1013 748 1017
rect 733 1012 737 1013
rect 664 1000 698 1004
rect 664 991 668 1000
rect 694 992 698 1000
rect 725 999 729 1004
rect 721 995 741 999
rect 656 979 660 983
rect 626 975 660 979
rect 676 976 680 980
rect 626 950 630 975
rect 639 965 643 969
rect 656 961 660 975
rect 618 938 622 942
rect 588 934 622 938
rect 638 935 642 939
rect 588 909 592 934
rect 601 924 605 928
rect 618 920 622 934
rect 580 897 584 901
rect 550 893 584 897
rect 600 894 604 898
rect 533 872 537 876
rect 550 868 554 893
rect 563 883 567 887
rect 580 879 584 893
rect 525 843 529 847
rect 542 839 546 860
rect 534 821 538 831
rect 572 821 576 871
rect 610 821 614 912
rect 648 821 652 953
rect 686 821 690 984
rect 706 977 710 981
rect 719 980 743 984
rect 725 975 729 980
rect 733 960 737 967
rect 764 960 768 1132
rect 788 1131 792 1132
rect 780 1118 784 1123
rect 776 1114 796 1118
rect 831 1113 835 1132
rect 854 1129 858 1132
rect 878 1126 882 1132
rect 873 1122 882 1126
rect 809 1108 813 1112
rect 809 1104 819 1108
rect 809 1092 813 1104
rect 827 1096 841 1100
rect 865 1098 873 1114
rect 878 1107 882 1122
rect 865 1094 921 1098
rect 865 1092 873 1094
rect 849 1088 873 1092
rect 834 1069 838 1080
rect 865 1074 873 1088
rect 917 1091 921 1094
rect 917 1087 944 1091
rect 794 1065 838 1069
rect 878 1066 882 1081
rect 917 1068 921 1087
rect 940 1084 944 1087
rect 964 1081 968 1087
rect 959 1077 968 1081
rect 794 1061 798 1065
rect 776 1054 780 1058
rect 818 1054 822 1060
rect 776 1050 785 1054
rect 813 1050 822 1054
rect 834 1055 838 1065
rect 873 1062 882 1066
rect 854 1055 858 1059
rect 878 1056 882 1062
rect 895 1063 899 1067
rect 895 1059 905 1063
rect 834 1051 858 1055
rect 776 1038 780 1050
rect 793 1042 805 1046
rect 794 1031 798 1042
rect 818 1036 822 1050
rect 895 1047 899 1059
rect 913 1051 927 1055
rect 951 1053 959 1069
rect 964 1062 968 1077
rect 987 1069 991 1289
rect 1297 1270 1301 1289
rect 1320 1286 1324 1289
rect 1344 1283 1348 1289
rect 1339 1279 1348 1283
rect 1275 1265 1279 1269
rect 1275 1261 1285 1265
rect 1275 1249 1279 1261
rect 1293 1253 1307 1257
rect 1331 1255 1339 1271
rect 1344 1264 1348 1279
rect 1356 1255 1360 1289
rect 1387 1270 1391 1289
rect 1410 1286 1414 1289
rect 1434 1283 1438 1289
rect 1429 1279 1438 1283
rect 1331 1251 1360 1255
rect 1365 1265 1369 1269
rect 1365 1261 1375 1265
rect 1331 1249 1339 1251
rect 1365 1249 1369 1261
rect 1383 1253 1397 1257
rect 1421 1255 1429 1271
rect 1434 1264 1438 1279
rect 1421 1251 1470 1255
rect 1421 1249 1429 1251
rect 1315 1245 1339 1249
rect 1405 1245 1429 1249
rect 999 1222 1200 1226
rect 999 1127 1003 1222
rect 1196 1221 1200 1222
rect 1196 1217 1223 1221
rect 1196 1198 1200 1217
rect 1219 1214 1223 1217
rect 1243 1211 1247 1217
rect 1238 1207 1247 1211
rect 1174 1193 1178 1197
rect 1174 1189 1184 1193
rect 1174 1177 1178 1189
rect 1192 1181 1206 1185
rect 1230 1180 1238 1199
rect 1243 1192 1247 1207
rect 1300 1212 1304 1237
rect 1331 1231 1339 1245
rect 1344 1223 1348 1238
rect 1339 1219 1348 1223
rect 1320 1212 1324 1216
rect 1344 1213 1348 1219
rect 1300 1208 1324 1212
rect 1390 1212 1394 1237
rect 1421 1231 1429 1245
rect 1434 1223 1438 1238
rect 1429 1219 1438 1223
rect 1410 1212 1414 1216
rect 1434 1213 1438 1219
rect 1390 1208 1414 1212
rect 1260 1200 1284 1204
rect 1266 1195 1270 1200
rect 1274 1180 1278 1187
rect 1300 1180 1304 1208
rect 1390 1199 1394 1208
rect 1390 1195 1454 1199
rect 1230 1177 1259 1180
rect 1214 1176 1259 1177
rect 1274 1176 1305 1180
rect 1214 1173 1238 1176
rect 1274 1175 1278 1176
rect 1007 1147 1031 1151
rect 1046 1147 1070 1151
rect 1086 1147 1110 1151
rect 1125 1147 1149 1151
rect 1166 1147 1190 1151
rect 1013 1142 1017 1147
rect 1052 1142 1056 1147
rect 1092 1142 1096 1147
rect 1131 1142 1135 1147
rect 1172 1142 1176 1147
rect 1021 1127 1025 1134
rect 1060 1127 1064 1134
rect 1100 1127 1104 1134
rect 1139 1127 1143 1134
rect 1180 1127 1184 1134
rect 1199 1140 1203 1165
rect 1230 1159 1238 1173
rect 1243 1151 1247 1166
rect 1266 1162 1270 1167
rect 1301 1163 1305 1176
rect 1262 1158 1282 1162
rect 1301 1159 1328 1163
rect 1360 1160 1418 1163
rect 1238 1147 1247 1151
rect 1219 1140 1223 1144
rect 1243 1141 1247 1147
rect 1199 1136 1223 1140
rect 1301 1140 1305 1159
rect 1324 1156 1328 1159
rect 1348 1153 1352 1159
rect 1343 1149 1352 1153
rect 1199 1127 1203 1136
rect 999 1123 1006 1127
rect 1021 1123 1045 1127
rect 1060 1123 1085 1127
rect 1100 1123 1124 1127
rect 1139 1123 1165 1127
rect 1180 1123 1203 1127
rect 1279 1135 1283 1139
rect 1279 1131 1289 1135
rect 1021 1122 1025 1123
rect 1060 1122 1064 1123
rect 1100 1122 1104 1123
rect 1139 1122 1143 1123
rect 1180 1122 1184 1123
rect 1279 1119 1283 1131
rect 1297 1123 1311 1127
rect 1335 1124 1343 1141
rect 1348 1134 1352 1149
rect 1360 1124 1364 1160
rect 1391 1159 1418 1160
rect 1391 1140 1395 1159
rect 1414 1156 1418 1159
rect 1438 1153 1442 1159
rect 1433 1149 1442 1153
rect 1335 1121 1364 1124
rect 1369 1135 1373 1139
rect 1369 1131 1379 1135
rect 1335 1119 1343 1121
rect 1369 1119 1373 1131
rect 1387 1123 1401 1127
rect 1425 1125 1433 1141
rect 1438 1134 1442 1149
rect 1450 1125 1454 1195
rect 1425 1121 1454 1125
rect 1425 1119 1433 1121
rect 1319 1115 1343 1119
rect 1409 1115 1433 1119
rect 1013 1109 1017 1114
rect 1052 1109 1056 1114
rect 1092 1109 1096 1114
rect 1131 1109 1135 1114
rect 1172 1109 1176 1114
rect 1009 1105 1029 1109
rect 1048 1105 1068 1109
rect 1088 1105 1108 1109
rect 1127 1105 1147 1109
rect 1168 1105 1188 1109
rect 995 1089 1019 1093
rect 1001 1084 1005 1089
rect 1009 1069 1013 1076
rect 1304 1082 1308 1107
rect 1335 1101 1343 1115
rect 1348 1093 1352 1108
rect 1343 1089 1352 1093
rect 1324 1082 1328 1086
rect 1348 1083 1352 1089
rect 1304 1078 1328 1082
rect 1394 1082 1398 1107
rect 1425 1101 1433 1115
rect 1438 1093 1442 1108
rect 1433 1089 1442 1093
rect 1414 1082 1418 1086
rect 1438 1083 1442 1089
rect 1394 1078 1418 1082
rect 1304 1069 1308 1078
rect 987 1065 994 1069
rect 1009 1065 1308 1069
rect 1394 1069 1398 1078
rect 1466 1069 1470 1251
rect 1394 1065 1470 1069
rect 1009 1064 1013 1065
rect 951 1049 971 1053
rect 1001 1051 1005 1056
rect 951 1047 959 1049
rect 997 1047 1017 1051
rect 935 1043 959 1047
rect 831 1037 858 1041
rect 831 1031 835 1037
rect 794 1027 835 1031
rect 854 1034 858 1037
rect 878 1031 882 1037
rect 873 1027 882 1031
rect 831 1018 835 1027
rect 809 1013 813 1017
rect 809 1009 819 1013
rect 809 997 813 1009
rect 827 1001 841 1005
rect 865 1003 873 1019
rect 878 1012 882 1027
rect 920 1010 924 1035
rect 951 1029 959 1043
rect 964 1021 968 1036
rect 959 1017 968 1021
rect 940 1010 944 1014
rect 964 1011 968 1017
rect 987 1033 1324 1037
rect 1356 1033 1414 1037
rect 920 1006 944 1010
rect 920 1003 924 1006
rect 865 999 924 1003
rect 865 997 873 999
rect 849 993 873 997
rect 834 960 838 985
rect 865 979 873 993
rect 878 971 882 986
rect 873 967 882 971
rect 854 960 858 964
rect 878 961 882 967
rect 712 956 718 960
rect 733 956 748 960
rect 764 956 858 960
rect 733 955 737 956
rect 725 942 729 947
rect 721 938 741 942
rect 719 923 743 927
rect 774 923 798 927
rect 725 918 729 923
rect 780 918 784 923
rect 733 903 737 910
rect 788 903 792 910
rect 712 899 718 903
rect 733 899 748 903
rect 764 899 773 903
rect 788 899 858 903
rect 733 898 737 899
rect 725 885 729 890
rect 721 881 741 885
rect 719 866 743 870
rect 725 861 729 866
rect 733 846 737 853
rect 712 842 718 846
rect 733 842 748 846
rect 733 841 737 842
rect 725 828 729 833
rect 721 824 741 828
rect 513 814 521 818
rect 534 817 690 821
rect 534 810 538 817
rect 405 799 461 803
rect 405 797 413 799
rect 389 793 413 797
rect 374 774 378 785
rect 405 779 413 793
rect 457 796 461 799
rect 526 796 530 802
rect 457 792 484 796
rect 522 792 542 796
rect 334 770 378 774
rect 418 771 422 786
rect 457 773 461 792
rect 480 789 484 792
rect 504 786 508 792
rect 499 782 508 786
rect 334 766 338 770
rect 316 759 320 763
rect 358 759 362 765
rect 316 755 325 759
rect 353 755 362 759
rect 374 760 378 770
rect 413 767 422 771
rect 394 760 398 764
rect 418 761 422 767
rect 435 768 439 772
rect 435 764 445 768
rect 374 756 398 760
rect 316 743 320 755
rect 333 747 345 751
rect 334 736 338 747
rect 358 741 362 755
rect 435 752 439 764
rect 453 756 467 760
rect 491 758 499 774
rect 504 767 508 782
rect 491 754 514 758
rect 491 752 499 754
rect 475 748 499 752
rect 371 742 398 746
rect 371 736 375 742
rect 334 732 375 736
rect 394 739 398 742
rect 418 736 422 742
rect 413 732 422 736
rect 371 723 375 732
rect 349 718 353 722
rect 349 714 359 718
rect 349 702 353 714
rect 367 706 381 710
rect 405 708 413 724
rect 418 717 422 732
rect 460 715 464 740
rect 491 734 499 748
rect 504 726 508 741
rect 499 722 508 726
rect 764 727 768 899
rect 788 898 792 899
rect 780 885 784 890
rect 776 881 796 885
rect 831 880 835 899
rect 854 896 858 899
rect 878 893 882 899
rect 873 889 882 893
rect 809 875 813 879
rect 809 871 819 875
rect 809 859 813 871
rect 827 863 841 867
rect 865 865 873 881
rect 878 874 882 889
rect 865 861 921 865
rect 865 859 873 861
rect 849 855 873 859
rect 834 836 838 847
rect 865 841 873 855
rect 917 858 921 861
rect 917 854 944 858
rect 794 832 838 836
rect 878 833 882 848
rect 917 835 921 854
rect 940 851 944 854
rect 964 848 968 854
rect 959 844 968 848
rect 794 828 798 832
rect 776 821 780 825
rect 818 821 822 827
rect 776 817 785 821
rect 813 817 822 821
rect 834 822 838 832
rect 873 829 882 833
rect 854 822 858 826
rect 878 823 882 829
rect 895 830 899 834
rect 895 826 905 830
rect 834 818 858 822
rect 776 805 780 817
rect 793 809 805 813
rect 794 798 798 809
rect 818 803 822 817
rect 895 814 899 826
rect 913 818 927 822
rect 951 820 959 836
rect 964 829 968 844
rect 951 816 971 820
rect 951 814 959 816
rect 935 810 959 814
rect 831 804 858 808
rect 831 798 835 804
rect 794 794 835 798
rect 854 801 858 804
rect 878 798 882 804
rect 873 794 882 798
rect 831 785 835 794
rect 809 780 813 784
rect 809 776 819 780
rect 809 764 813 776
rect 827 768 841 772
rect 865 770 873 786
rect 878 779 882 794
rect 920 777 924 802
rect 951 796 959 810
rect 987 813 991 1033
rect 1297 1014 1301 1033
rect 1320 1030 1324 1033
rect 1344 1027 1348 1033
rect 1339 1023 1348 1027
rect 1275 1009 1279 1013
rect 1275 1005 1285 1009
rect 1275 993 1279 1005
rect 1293 997 1307 1001
rect 1331 999 1339 1015
rect 1344 1008 1348 1023
rect 1356 999 1360 1033
rect 1387 1014 1391 1033
rect 1410 1030 1414 1033
rect 1434 1027 1438 1033
rect 1429 1023 1438 1027
rect 1331 995 1360 999
rect 1365 1009 1369 1013
rect 1365 1005 1375 1009
rect 1331 993 1339 995
rect 1365 993 1369 1005
rect 1383 997 1397 1001
rect 1421 999 1429 1015
rect 1434 1008 1438 1023
rect 1421 995 1470 999
rect 1421 993 1429 995
rect 1315 989 1339 993
rect 1405 989 1429 993
rect 999 966 1200 970
rect 999 871 1003 966
rect 1196 965 1200 966
rect 1196 961 1223 965
rect 1196 942 1200 961
rect 1219 958 1223 961
rect 1243 955 1247 961
rect 1238 951 1247 955
rect 1174 937 1178 941
rect 1174 933 1184 937
rect 1174 921 1178 933
rect 1192 925 1206 929
rect 1230 924 1238 943
rect 1243 936 1247 951
rect 1300 956 1304 981
rect 1331 975 1339 989
rect 1344 967 1348 982
rect 1339 963 1348 967
rect 1320 956 1324 960
rect 1344 957 1348 963
rect 1300 952 1324 956
rect 1390 956 1394 981
rect 1421 975 1429 989
rect 1434 967 1438 982
rect 1429 963 1438 967
rect 1410 956 1414 960
rect 1434 957 1438 963
rect 1390 952 1414 956
rect 1260 944 1284 948
rect 1266 939 1270 944
rect 1274 924 1278 931
rect 1300 924 1304 952
rect 1390 943 1394 952
rect 1390 939 1454 943
rect 1230 921 1259 924
rect 1214 920 1259 921
rect 1274 920 1305 924
rect 1214 917 1238 920
rect 1274 919 1278 920
rect 1007 891 1031 895
rect 1046 891 1070 895
rect 1086 891 1110 895
rect 1125 891 1149 895
rect 1166 891 1190 895
rect 1013 886 1017 891
rect 1052 886 1056 891
rect 1092 886 1096 891
rect 1131 886 1135 891
rect 1172 886 1176 891
rect 1021 871 1025 878
rect 1060 871 1064 878
rect 1100 871 1104 878
rect 1139 871 1143 878
rect 1180 871 1184 878
rect 1199 884 1203 909
rect 1230 903 1238 917
rect 1243 895 1247 910
rect 1266 906 1270 911
rect 1301 907 1305 920
rect 1262 902 1282 906
rect 1301 903 1328 907
rect 1360 904 1418 907
rect 1238 891 1247 895
rect 1219 884 1223 888
rect 1243 885 1247 891
rect 1199 880 1223 884
rect 1301 884 1305 903
rect 1324 900 1328 903
rect 1348 897 1352 903
rect 1343 893 1352 897
rect 1199 871 1203 880
rect 999 867 1006 871
rect 1021 867 1045 871
rect 1060 867 1085 871
rect 1100 867 1124 871
rect 1139 867 1165 871
rect 1180 867 1203 871
rect 1279 879 1283 883
rect 1279 875 1289 879
rect 1021 866 1025 867
rect 1060 866 1064 867
rect 1100 866 1104 867
rect 1139 866 1143 867
rect 1180 866 1184 867
rect 1279 863 1283 875
rect 1297 867 1311 871
rect 1335 868 1343 885
rect 1348 878 1352 893
rect 1360 868 1364 904
rect 1391 903 1418 904
rect 1391 884 1395 903
rect 1414 900 1418 903
rect 1438 897 1442 903
rect 1433 893 1442 897
rect 1335 865 1364 868
rect 1369 879 1373 883
rect 1369 875 1379 879
rect 1335 863 1343 865
rect 1369 863 1373 875
rect 1387 867 1401 871
rect 1425 869 1433 885
rect 1438 878 1442 893
rect 1450 869 1454 939
rect 1425 865 1454 869
rect 1425 863 1433 865
rect 1319 859 1343 863
rect 1409 859 1433 863
rect 1013 853 1017 858
rect 1052 853 1056 858
rect 1092 853 1096 858
rect 1131 853 1135 858
rect 1172 853 1176 858
rect 1009 849 1029 853
rect 1048 849 1068 853
rect 1088 849 1108 853
rect 1127 849 1147 853
rect 1168 849 1188 853
rect 995 833 1019 837
rect 1001 828 1005 833
rect 1009 813 1013 820
rect 1304 826 1308 851
rect 1335 845 1343 859
rect 1348 837 1352 852
rect 1343 833 1352 837
rect 1324 826 1328 830
rect 1348 827 1352 833
rect 1304 822 1328 826
rect 1394 826 1398 851
rect 1425 845 1433 859
rect 1438 837 1442 852
rect 1433 833 1442 837
rect 1414 826 1418 830
rect 1438 827 1442 833
rect 1394 822 1418 826
rect 1304 813 1308 822
rect 987 809 994 813
rect 1009 809 1308 813
rect 1394 813 1398 822
rect 1466 813 1470 995
rect 1394 809 1470 813
rect 1009 808 1013 809
rect 964 788 968 803
rect 1001 795 1005 800
rect 997 791 1017 795
rect 959 784 968 788
rect 940 777 944 781
rect 964 778 968 784
rect 920 773 944 777
rect 987 777 1324 781
rect 1356 777 1414 781
rect 920 770 924 773
rect 865 766 924 770
rect 865 764 873 766
rect 849 760 873 764
rect 834 727 838 752
rect 865 746 873 760
rect 878 738 882 753
rect 873 734 882 738
rect 854 727 858 731
rect 878 728 882 734
rect 764 723 858 727
rect 480 715 484 719
rect 504 716 508 722
rect 460 711 484 715
rect 460 708 464 711
rect 405 704 464 708
rect 405 702 413 704
rect 389 698 413 702
rect 374 665 378 690
rect 405 684 413 698
rect 418 676 422 691
rect 774 690 798 694
rect 780 685 784 690
rect 413 672 422 676
rect 394 665 398 669
rect 418 666 422 672
rect 788 670 792 677
rect 764 666 773 670
rect 788 666 858 670
rect 304 661 398 665
rect 212 652 288 656
rect -173 651 -169 652
rect -181 638 -177 643
rect -185 634 -165 638
rect 326 629 353 633
rect -195 620 142 624
rect 174 620 232 624
rect -195 400 -191 620
rect 115 601 119 620
rect 138 617 142 620
rect 162 614 166 620
rect 157 610 166 614
rect 93 596 97 600
rect 93 592 103 596
rect 93 580 97 592
rect 111 584 125 588
rect 149 586 157 602
rect 162 595 166 610
rect 174 586 178 620
rect 205 601 209 620
rect 228 617 232 620
rect 252 614 256 620
rect 247 610 256 614
rect 149 582 178 586
rect 183 596 187 600
rect 183 592 193 596
rect 149 580 157 582
rect 183 580 187 592
rect 201 584 215 588
rect 239 586 247 602
rect 252 595 256 610
rect 326 610 330 629
rect 349 626 353 629
rect 373 623 377 629
rect 368 619 377 623
rect 304 605 308 609
rect 304 601 314 605
rect 304 589 308 601
rect 322 593 336 597
rect 360 595 368 611
rect 373 604 377 619
rect 391 615 415 619
rect 397 610 401 615
rect 405 595 409 602
rect 360 591 390 595
rect 405 591 426 595
rect 360 589 368 591
rect 405 590 409 591
rect 239 582 288 586
rect 344 585 368 589
rect 239 580 247 582
rect 133 576 157 580
rect 223 576 247 580
rect -183 553 18 557
rect -183 458 -179 553
rect 14 552 18 553
rect 14 548 41 552
rect 14 529 18 548
rect 37 545 41 548
rect 61 542 65 548
rect 56 538 65 542
rect -8 524 -4 528
rect -8 520 2 524
rect -8 508 -4 520
rect 10 512 24 516
rect 48 511 56 530
rect 61 523 65 538
rect 118 543 122 568
rect 149 562 157 576
rect 162 554 166 569
rect 157 550 166 554
rect 138 543 142 547
rect 162 544 166 550
rect 118 539 142 543
rect 208 543 212 568
rect 239 562 247 576
rect 252 554 256 569
rect 247 550 256 554
rect 228 543 232 547
rect 252 544 256 550
rect 208 539 232 543
rect 78 531 102 535
rect 84 526 88 531
rect 92 511 96 518
rect 118 511 122 539
rect 208 530 212 539
rect 208 526 272 530
rect 48 508 77 511
rect 32 507 77 508
rect 92 507 123 511
rect 32 504 56 507
rect 92 506 96 507
rect -175 478 -151 482
rect -136 478 -112 482
rect -96 478 -72 482
rect -57 478 -33 482
rect -16 478 8 482
rect -169 473 -165 478
rect -130 473 -126 478
rect -90 473 -86 478
rect -51 473 -47 478
rect -10 473 -6 478
rect -161 458 -157 465
rect -122 458 -118 465
rect -82 458 -78 465
rect -43 458 -39 465
rect -2 458 2 465
rect 17 471 21 496
rect 48 490 56 504
rect 61 482 65 497
rect 84 493 88 498
rect 119 494 123 507
rect 80 489 100 493
rect 119 490 146 494
rect 178 491 236 494
rect 56 478 65 482
rect 37 471 41 475
rect 61 472 65 478
rect 17 467 41 471
rect 119 471 123 490
rect 142 487 146 490
rect 166 484 170 490
rect 161 480 170 484
rect 17 458 21 467
rect -183 454 -176 458
rect -161 454 -137 458
rect -122 454 -97 458
rect -82 454 -58 458
rect -43 454 -17 458
rect -2 454 21 458
rect 97 466 101 470
rect 97 462 107 466
rect -161 453 -157 454
rect -122 453 -118 454
rect -82 453 -78 454
rect -43 453 -39 454
rect -2 453 2 454
rect 97 450 101 462
rect 115 454 129 458
rect 153 455 161 472
rect 166 465 170 480
rect 178 455 182 491
rect 209 490 236 491
rect 209 471 213 490
rect 232 487 236 490
rect 256 484 260 490
rect 251 480 260 484
rect 153 452 182 455
rect 187 466 191 470
rect 187 462 197 466
rect 153 450 161 452
rect 187 450 191 462
rect 205 454 219 458
rect 243 456 251 472
rect 256 465 260 480
rect 268 456 272 526
rect 243 452 272 456
rect 243 450 251 452
rect 137 446 161 450
rect 227 446 251 450
rect -169 440 -165 445
rect -130 440 -126 445
rect -90 440 -86 445
rect -51 440 -47 445
rect -10 440 -6 445
rect -173 436 -153 440
rect -134 436 -114 440
rect -94 436 -74 440
rect -55 436 -35 440
rect -14 436 6 440
rect -187 420 -163 424
rect -181 415 -177 420
rect -173 400 -169 407
rect 122 413 126 438
rect 153 432 161 446
rect 166 424 170 439
rect 161 420 170 424
rect 142 413 146 417
rect 166 414 170 420
rect 122 409 146 413
rect 212 413 216 438
rect 243 432 251 446
rect 256 424 260 439
rect 251 420 260 424
rect 232 413 236 417
rect 256 414 260 420
rect 212 409 236 413
rect 122 400 126 409
rect -195 396 -188 400
rect -173 396 126 400
rect 212 400 216 409
rect 284 400 288 582
rect 329 552 333 577
rect 360 571 368 585
rect 373 563 377 578
rect 397 577 401 582
rect 393 573 413 577
rect 368 559 377 563
rect 349 552 353 556
rect 373 553 377 559
rect 329 548 353 552
rect 314 526 338 530
rect 320 521 324 526
rect 328 506 332 513
rect 212 396 288 400
rect 304 502 313 506
rect 328 502 398 506
rect -173 395 -169 396
rect -181 382 -177 387
rect -185 378 -165 382
rect -195 364 142 368
rect 174 364 232 368
rect -195 144 -191 364
rect 115 345 119 364
rect 138 361 142 364
rect 162 358 166 364
rect 157 354 166 358
rect 93 340 97 344
rect 93 336 103 340
rect 93 324 97 336
rect 111 328 125 332
rect 149 330 157 346
rect 162 339 166 354
rect 174 330 178 364
rect 205 345 209 364
rect 228 361 232 364
rect 252 358 256 364
rect 247 354 256 358
rect 149 326 178 330
rect 183 340 187 344
rect 183 336 193 340
rect 149 324 157 326
rect 183 324 187 336
rect 201 328 215 332
rect 239 330 247 346
rect 252 339 256 354
rect 304 330 308 502
rect 328 501 332 502
rect 320 488 324 493
rect 316 484 336 488
rect 371 483 375 502
rect 394 499 398 502
rect 418 496 422 502
rect 413 492 422 496
rect 349 478 353 482
rect 349 474 359 478
rect 349 462 353 474
rect 367 466 381 470
rect 405 468 413 484
rect 418 477 422 492
rect 764 494 768 666
rect 788 665 792 666
rect 780 652 784 657
rect 776 648 796 652
rect 831 647 835 666
rect 854 663 858 666
rect 878 660 882 666
rect 873 656 882 660
rect 809 642 813 646
rect 809 638 819 642
rect 809 626 813 638
rect 827 630 841 634
rect 865 632 873 648
rect 878 641 882 656
rect 865 628 921 632
rect 865 626 873 628
rect 849 622 873 626
rect 834 603 838 614
rect 865 608 873 622
rect 917 625 921 628
rect 917 621 944 625
rect 794 599 838 603
rect 878 600 882 615
rect 917 602 921 621
rect 940 618 944 621
rect 964 615 968 621
rect 959 611 968 615
rect 794 595 798 599
rect 776 588 780 592
rect 818 588 822 594
rect 776 584 785 588
rect 813 584 822 588
rect 834 589 838 599
rect 873 596 882 600
rect 854 589 858 593
rect 878 590 882 596
rect 895 597 899 601
rect 895 593 905 597
rect 834 585 858 589
rect 776 572 780 584
rect 793 576 805 580
rect 794 565 798 576
rect 818 570 822 584
rect 895 581 899 593
rect 913 585 927 589
rect 951 587 959 603
rect 964 596 968 611
rect 951 583 971 587
rect 951 581 959 583
rect 935 577 959 581
rect 831 571 858 575
rect 831 565 835 571
rect 794 561 835 565
rect 854 568 858 571
rect 878 565 882 571
rect 873 561 882 565
rect 831 552 835 561
rect 809 547 813 551
rect 809 543 819 547
rect 809 531 813 543
rect 827 535 841 539
rect 865 537 873 553
rect 878 546 882 561
rect 920 544 924 569
rect 951 563 959 577
rect 964 555 968 570
rect 959 551 968 555
rect 987 557 991 777
rect 1297 758 1301 777
rect 1320 774 1324 777
rect 1344 771 1348 777
rect 1339 767 1348 771
rect 1275 753 1279 757
rect 1275 749 1285 753
rect 1275 737 1279 749
rect 1293 741 1307 745
rect 1331 743 1339 759
rect 1344 752 1348 767
rect 1356 743 1360 777
rect 1387 758 1391 777
rect 1410 774 1414 777
rect 1434 771 1438 777
rect 1429 767 1438 771
rect 1331 739 1360 743
rect 1365 753 1369 757
rect 1365 749 1375 753
rect 1331 737 1339 739
rect 1365 737 1369 749
rect 1383 741 1397 745
rect 1421 743 1429 759
rect 1434 752 1438 767
rect 1421 739 1470 743
rect 1421 737 1429 739
rect 1315 733 1339 737
rect 1405 733 1429 737
rect 999 710 1200 714
rect 999 615 1003 710
rect 1196 709 1200 710
rect 1196 705 1223 709
rect 1196 686 1200 705
rect 1219 702 1223 705
rect 1243 699 1247 705
rect 1238 695 1247 699
rect 1174 681 1178 685
rect 1174 677 1184 681
rect 1174 665 1178 677
rect 1192 669 1206 673
rect 1230 668 1238 687
rect 1243 680 1247 695
rect 1300 700 1304 725
rect 1331 719 1339 733
rect 1344 711 1348 726
rect 1339 707 1348 711
rect 1320 700 1324 704
rect 1344 701 1348 707
rect 1300 696 1324 700
rect 1390 700 1394 725
rect 1421 719 1429 733
rect 1434 711 1438 726
rect 1429 707 1438 711
rect 1410 700 1414 704
rect 1434 701 1438 707
rect 1390 696 1414 700
rect 1260 688 1284 692
rect 1266 683 1270 688
rect 1274 668 1278 675
rect 1300 668 1304 696
rect 1390 687 1394 696
rect 1390 683 1454 687
rect 1230 665 1259 668
rect 1214 664 1259 665
rect 1274 664 1305 668
rect 1214 661 1238 664
rect 1274 663 1278 664
rect 1007 635 1031 639
rect 1046 635 1070 639
rect 1086 635 1110 639
rect 1125 635 1149 639
rect 1166 635 1190 639
rect 1013 630 1017 635
rect 1052 630 1056 635
rect 1092 630 1096 635
rect 1131 630 1135 635
rect 1172 630 1176 635
rect 1021 615 1025 622
rect 1060 615 1064 622
rect 1100 615 1104 622
rect 1139 615 1143 622
rect 1180 615 1184 622
rect 1199 628 1203 653
rect 1230 647 1238 661
rect 1243 639 1247 654
rect 1266 650 1270 655
rect 1301 651 1305 664
rect 1262 646 1282 650
rect 1301 647 1328 651
rect 1360 648 1418 651
rect 1238 635 1247 639
rect 1219 628 1223 632
rect 1243 629 1247 635
rect 1199 624 1223 628
rect 1301 628 1305 647
rect 1324 644 1328 647
rect 1348 641 1352 647
rect 1343 637 1352 641
rect 1199 615 1203 624
rect 999 611 1006 615
rect 1021 611 1045 615
rect 1060 611 1085 615
rect 1100 611 1124 615
rect 1139 611 1165 615
rect 1180 611 1203 615
rect 1279 623 1283 627
rect 1279 619 1289 623
rect 1021 610 1025 611
rect 1060 610 1064 611
rect 1100 610 1104 611
rect 1139 610 1143 611
rect 1180 610 1184 611
rect 1279 607 1283 619
rect 1297 611 1311 615
rect 1335 612 1343 629
rect 1348 622 1352 637
rect 1360 612 1364 648
rect 1391 647 1418 648
rect 1391 628 1395 647
rect 1414 644 1418 647
rect 1438 641 1442 647
rect 1433 637 1442 641
rect 1335 609 1364 612
rect 1369 623 1373 627
rect 1369 619 1379 623
rect 1335 607 1343 609
rect 1369 607 1373 619
rect 1387 611 1401 615
rect 1425 613 1433 629
rect 1438 622 1442 637
rect 1450 613 1454 683
rect 1425 609 1454 613
rect 1425 607 1433 609
rect 1319 603 1343 607
rect 1409 603 1433 607
rect 1013 597 1017 602
rect 1052 597 1056 602
rect 1092 597 1096 602
rect 1131 597 1135 602
rect 1172 597 1176 602
rect 1009 593 1029 597
rect 1048 593 1068 597
rect 1088 593 1108 597
rect 1127 593 1147 597
rect 1168 593 1188 597
rect 995 577 1019 581
rect 1001 572 1005 577
rect 1009 557 1013 564
rect 1304 570 1308 595
rect 1335 589 1343 603
rect 1348 581 1352 596
rect 1343 577 1352 581
rect 1324 570 1328 574
rect 1348 571 1352 577
rect 1304 566 1328 570
rect 1394 570 1398 595
rect 1425 589 1433 603
rect 1438 581 1442 596
rect 1433 577 1442 581
rect 1414 570 1418 574
rect 1438 571 1442 577
rect 1394 566 1418 570
rect 1304 557 1308 566
rect 987 553 994 557
rect 1009 553 1308 557
rect 1394 557 1398 566
rect 1466 557 1470 739
rect 1394 553 1470 557
rect 1009 552 1013 553
rect 940 544 944 548
rect 964 545 968 551
rect 920 540 944 544
rect 920 537 924 540
rect 1001 539 1005 544
rect 865 533 924 537
rect 997 535 1017 539
rect 865 531 873 533
rect 849 527 873 531
rect 774 514 798 518
rect 780 509 784 514
rect 788 494 792 501
rect 834 494 838 519
rect 865 513 873 527
rect 987 521 1324 525
rect 1356 521 1414 525
rect 878 505 882 520
rect 873 501 882 505
rect 854 494 858 498
rect 878 495 882 501
rect 764 490 773 494
rect 788 490 858 494
rect 788 489 792 490
rect 780 476 784 481
rect 776 472 796 476
rect 405 464 461 468
rect 405 462 413 464
rect 389 458 413 462
rect 374 439 378 450
rect 405 444 413 458
rect 457 461 461 464
rect 457 457 484 461
rect 334 435 378 439
rect 418 436 422 451
rect 457 438 461 457
rect 480 454 484 457
rect 504 451 508 457
rect 499 447 508 451
rect 334 431 338 435
rect 316 424 320 428
rect 358 424 362 430
rect 316 420 325 424
rect 353 420 362 424
rect 374 425 378 435
rect 413 432 422 436
rect 394 425 398 429
rect 418 426 422 432
rect 435 433 439 437
rect 435 429 445 433
rect 374 421 398 425
rect 316 408 320 420
rect 333 412 345 416
rect 334 401 338 412
rect 358 406 362 420
rect 435 417 439 429
rect 453 421 467 425
rect 491 423 499 439
rect 504 432 508 447
rect 491 419 514 423
rect 491 417 499 419
rect 475 413 499 417
rect 371 407 398 411
rect 371 401 375 407
rect 334 397 375 401
rect 394 404 398 407
rect 418 401 422 407
rect 413 397 422 401
rect 371 388 375 397
rect 349 383 353 387
rect 349 379 359 383
rect 349 367 353 379
rect 367 371 381 375
rect 405 373 413 389
rect 418 382 422 397
rect 460 380 464 405
rect 491 399 499 413
rect 504 391 508 406
rect 499 387 508 391
rect 480 380 484 384
rect 504 381 508 387
rect 460 376 484 380
rect 460 373 464 376
rect 405 369 464 373
rect 405 367 413 369
rect 389 363 413 367
rect 374 330 378 355
rect 405 349 413 363
rect 418 341 422 356
rect 413 337 422 341
rect 394 330 398 334
rect 418 331 422 337
rect 239 326 288 330
rect 304 326 398 330
rect 239 324 247 326
rect 133 320 157 324
rect 223 320 247 324
rect -183 297 18 301
rect -183 202 -179 297
rect 14 296 18 297
rect 14 292 41 296
rect 14 273 18 292
rect 37 289 41 292
rect 61 286 65 292
rect 56 282 65 286
rect -8 268 -4 272
rect -8 264 2 268
rect -8 252 -4 264
rect 10 256 24 260
rect 48 255 56 274
rect 61 267 65 282
rect 118 287 122 312
rect 149 306 157 320
rect 162 298 166 313
rect 157 294 166 298
rect 138 287 142 291
rect 162 288 166 294
rect 118 283 142 287
rect 208 287 212 312
rect 239 306 247 320
rect 252 298 256 313
rect 247 294 256 298
rect 228 287 232 291
rect 252 288 256 294
rect 208 283 232 287
rect 78 275 102 279
rect 84 270 88 275
rect 92 255 96 262
rect 118 255 122 283
rect 208 274 212 283
rect 208 270 272 274
rect 48 252 77 255
rect 32 251 77 252
rect 92 251 123 255
rect 32 248 56 251
rect 92 250 96 251
rect -175 222 -151 226
rect -136 222 -112 226
rect -96 222 -72 226
rect -57 222 -33 226
rect -16 222 8 226
rect -169 217 -165 222
rect -130 217 -126 222
rect -90 217 -86 222
rect -51 217 -47 222
rect -10 217 -6 222
rect -161 202 -157 209
rect -122 202 -118 209
rect -82 202 -78 209
rect -43 202 -39 209
rect -2 202 2 209
rect 17 215 21 240
rect 48 234 56 248
rect 61 226 65 241
rect 84 237 88 242
rect 119 238 123 251
rect 80 233 100 237
rect 119 234 146 238
rect 178 235 236 238
rect 56 222 65 226
rect 37 215 41 219
rect 61 216 65 222
rect 17 211 41 215
rect 119 215 123 234
rect 142 231 146 234
rect 166 228 170 234
rect 161 224 170 228
rect 17 202 21 211
rect -183 198 -176 202
rect -161 198 -137 202
rect -122 198 -97 202
rect -82 198 -58 202
rect -43 198 -17 202
rect -2 198 21 202
rect 97 210 101 214
rect 97 206 107 210
rect -161 197 -157 198
rect -122 197 -118 198
rect -82 197 -78 198
rect -43 197 -39 198
rect -2 197 2 198
rect 97 194 101 206
rect 115 198 129 202
rect 153 199 161 216
rect 166 209 170 224
rect 178 199 182 235
rect 209 234 236 235
rect 209 215 213 234
rect 232 231 236 234
rect 256 228 260 234
rect 251 224 260 228
rect 153 196 182 199
rect 187 210 191 214
rect 187 206 197 210
rect 153 194 161 196
rect 187 194 191 206
rect 205 198 219 202
rect 243 200 251 216
rect 256 209 260 224
rect 268 200 272 270
rect 243 196 272 200
rect 243 194 251 196
rect 137 190 161 194
rect 227 190 251 194
rect -169 184 -165 189
rect -130 184 -126 189
rect -90 184 -86 189
rect -51 184 -47 189
rect -10 184 -6 189
rect -173 180 -153 184
rect -134 180 -114 184
rect -94 180 -74 184
rect -55 180 -35 184
rect -14 180 6 184
rect -187 164 -163 168
rect -181 159 -177 164
rect -173 144 -169 151
rect 122 157 126 182
rect 153 176 161 190
rect 166 168 170 183
rect 161 164 170 168
rect 142 157 146 161
rect 166 158 170 164
rect 122 153 146 157
rect 212 157 216 182
rect 243 176 251 190
rect 256 168 260 183
rect 251 164 260 168
rect 232 157 236 161
rect 256 158 260 164
rect 212 153 236 157
rect 122 144 126 153
rect -195 140 -188 144
rect -173 140 126 144
rect 212 144 216 153
rect 284 144 288 326
rect 987 301 991 521
rect 1297 502 1301 521
rect 1320 518 1324 521
rect 1344 515 1348 521
rect 1339 511 1348 515
rect 1275 497 1279 501
rect 1275 493 1285 497
rect 1275 481 1279 493
rect 1293 485 1307 489
rect 1331 487 1339 503
rect 1344 496 1348 511
rect 1356 487 1360 521
rect 1387 502 1391 521
rect 1410 518 1414 521
rect 1434 515 1438 521
rect 1429 511 1438 515
rect 1331 483 1360 487
rect 1365 497 1369 501
rect 1365 493 1375 497
rect 1331 481 1339 483
rect 1365 481 1369 493
rect 1383 485 1397 489
rect 1421 487 1429 503
rect 1434 496 1438 511
rect 1421 483 1470 487
rect 1421 481 1429 483
rect 1315 477 1339 481
rect 1405 477 1429 481
rect 999 454 1200 458
rect 999 359 1003 454
rect 1196 453 1200 454
rect 1196 449 1223 453
rect 1196 430 1200 449
rect 1219 446 1223 449
rect 1243 443 1247 449
rect 1238 439 1247 443
rect 1174 425 1178 429
rect 1174 421 1184 425
rect 1174 409 1178 421
rect 1192 413 1206 417
rect 1230 412 1238 431
rect 1243 424 1247 439
rect 1300 444 1304 469
rect 1331 463 1339 477
rect 1344 455 1348 470
rect 1339 451 1348 455
rect 1320 444 1324 448
rect 1344 445 1348 451
rect 1300 440 1324 444
rect 1390 444 1394 469
rect 1421 463 1429 477
rect 1434 455 1438 470
rect 1429 451 1438 455
rect 1410 444 1414 448
rect 1434 445 1438 451
rect 1390 440 1414 444
rect 1260 432 1284 436
rect 1266 427 1270 432
rect 1274 412 1278 419
rect 1300 412 1304 440
rect 1390 431 1394 440
rect 1390 427 1454 431
rect 1230 409 1259 412
rect 1214 408 1259 409
rect 1274 408 1305 412
rect 1214 405 1238 408
rect 1274 407 1278 408
rect 1007 379 1031 383
rect 1046 379 1070 383
rect 1086 379 1110 383
rect 1125 379 1149 383
rect 1166 379 1190 383
rect 1013 374 1017 379
rect 1052 374 1056 379
rect 1092 374 1096 379
rect 1131 374 1135 379
rect 1172 374 1176 379
rect 1021 359 1025 366
rect 1060 359 1064 366
rect 1100 359 1104 366
rect 1139 359 1143 366
rect 1180 359 1184 366
rect 1199 372 1203 397
rect 1230 391 1238 405
rect 1243 383 1247 398
rect 1266 394 1270 399
rect 1301 395 1305 408
rect 1262 390 1282 394
rect 1301 391 1328 395
rect 1360 392 1418 395
rect 1238 379 1247 383
rect 1219 372 1223 376
rect 1243 373 1247 379
rect 1199 368 1223 372
rect 1301 372 1305 391
rect 1324 388 1328 391
rect 1348 385 1352 391
rect 1343 381 1352 385
rect 1199 359 1203 368
rect 999 355 1006 359
rect 1021 355 1045 359
rect 1060 355 1085 359
rect 1100 355 1124 359
rect 1139 355 1165 359
rect 1180 355 1203 359
rect 1279 367 1283 371
rect 1279 363 1289 367
rect 1021 354 1025 355
rect 1060 354 1064 355
rect 1100 354 1104 355
rect 1139 354 1143 355
rect 1180 354 1184 355
rect 1279 351 1283 363
rect 1297 355 1311 359
rect 1335 356 1343 373
rect 1348 366 1352 381
rect 1360 356 1364 392
rect 1391 391 1418 392
rect 1391 372 1395 391
rect 1414 388 1418 391
rect 1438 385 1442 391
rect 1433 381 1442 385
rect 1335 353 1364 356
rect 1369 367 1373 371
rect 1369 363 1379 367
rect 1335 351 1343 353
rect 1369 351 1373 363
rect 1387 355 1401 359
rect 1425 357 1433 373
rect 1438 366 1442 381
rect 1450 357 1454 427
rect 1425 353 1454 357
rect 1425 351 1433 353
rect 1319 347 1343 351
rect 1409 347 1433 351
rect 1013 341 1017 346
rect 1052 341 1056 346
rect 1092 341 1096 346
rect 1131 341 1135 346
rect 1172 341 1176 346
rect 1009 337 1029 341
rect 1048 337 1068 341
rect 1088 337 1108 341
rect 1127 337 1147 341
rect 1168 337 1188 341
rect 995 321 1019 325
rect 1001 316 1005 321
rect 1009 301 1013 308
rect 1304 314 1308 339
rect 1335 333 1343 347
rect 1348 325 1352 340
rect 1343 321 1352 325
rect 1324 314 1328 318
rect 1348 315 1352 321
rect 1304 310 1328 314
rect 1394 314 1398 339
rect 1425 333 1433 347
rect 1438 325 1442 340
rect 1433 321 1442 325
rect 1414 314 1418 318
rect 1438 315 1442 321
rect 1394 310 1418 314
rect 1304 301 1308 310
rect 326 294 353 298
rect 987 297 994 301
rect 1009 297 1308 301
rect 1394 301 1398 310
rect 1466 301 1470 483
rect 1394 297 1470 301
rect 1009 296 1013 297
rect 326 275 330 294
rect 349 291 353 294
rect 373 288 377 294
rect 368 284 377 288
rect 304 270 308 274
rect 304 266 314 270
rect 304 254 308 266
rect 322 258 336 262
rect 360 260 368 276
rect 373 269 377 284
rect 391 280 415 284
rect 1001 283 1005 288
rect 397 275 401 280
rect 997 279 1017 283
rect 405 260 409 267
rect 360 256 390 260
rect 405 256 426 260
rect 360 254 368 256
rect 405 255 409 256
rect 344 250 368 254
rect 329 217 333 242
rect 360 236 368 250
rect 373 228 377 243
rect 397 242 401 247
rect 393 238 413 242
rect 368 224 377 228
rect 349 217 353 221
rect 373 218 377 224
rect 329 213 353 217
rect 212 140 288 144
rect -173 139 -169 140
rect -181 126 -177 131
rect -185 122 -165 126
rect -195 108 142 112
rect 174 108 232 112
rect -195 -112 -191 108
rect 115 89 119 108
rect 138 105 142 108
rect 162 102 166 108
rect 157 98 166 102
rect 93 84 97 88
rect 93 80 103 84
rect 93 68 97 80
rect 111 72 125 76
rect 149 74 157 90
rect 162 83 166 98
rect 174 74 178 108
rect 205 89 209 108
rect 228 105 232 108
rect 252 102 256 108
rect 247 98 256 102
rect 149 70 178 74
rect 183 84 187 88
rect 183 80 193 84
rect 149 68 157 70
rect 183 68 187 80
rect 201 72 215 76
rect 239 74 247 90
rect 252 83 256 98
rect 239 70 288 74
rect 239 68 247 70
rect 133 64 157 68
rect 223 64 247 68
rect -183 41 18 45
rect -183 -54 -179 41
rect 14 40 18 41
rect 14 36 41 40
rect 14 17 18 36
rect 37 33 41 36
rect 61 30 65 36
rect 56 26 65 30
rect -8 12 -4 16
rect -8 8 2 12
rect -8 -4 -4 8
rect 10 0 24 4
rect 48 -1 56 18
rect 61 11 65 26
rect 118 31 122 56
rect 149 50 157 64
rect 162 42 166 57
rect 157 38 166 42
rect 138 31 142 35
rect 162 32 166 38
rect 118 27 142 31
rect 208 31 212 56
rect 239 50 247 64
rect 252 42 256 57
rect 247 38 256 42
rect 228 31 232 35
rect 252 32 256 38
rect 208 27 232 31
rect 78 19 102 23
rect 84 14 88 19
rect 92 -1 96 6
rect 118 -1 122 27
rect 208 18 212 27
rect 208 14 272 18
rect 48 -4 77 -1
rect 32 -5 77 -4
rect 92 -5 123 -1
rect 32 -8 56 -5
rect 92 -6 96 -5
rect -175 -34 -151 -30
rect -136 -34 -112 -30
rect -96 -34 -72 -30
rect -57 -34 -33 -30
rect -16 -34 8 -30
rect -169 -39 -165 -34
rect -130 -39 -126 -34
rect -90 -39 -86 -34
rect -51 -39 -47 -34
rect -10 -39 -6 -34
rect -161 -54 -157 -47
rect -122 -54 -118 -47
rect -82 -54 -78 -47
rect -43 -54 -39 -47
rect -2 -54 2 -47
rect 17 -41 21 -16
rect 48 -22 56 -8
rect 61 -30 65 -15
rect 84 -19 88 -14
rect 119 -18 123 -5
rect 80 -23 100 -19
rect 119 -22 146 -18
rect 178 -21 236 -18
rect 56 -34 65 -30
rect 37 -41 41 -37
rect 61 -40 65 -34
rect 17 -45 41 -41
rect 119 -41 123 -22
rect 142 -25 146 -22
rect 166 -28 170 -22
rect 161 -32 170 -28
rect 17 -54 21 -45
rect -183 -58 -176 -54
rect -161 -58 -137 -54
rect -122 -58 -97 -54
rect -82 -58 -58 -54
rect -43 -58 -17 -54
rect -2 -58 21 -54
rect 97 -46 101 -42
rect 97 -50 107 -46
rect -161 -59 -157 -58
rect -122 -59 -118 -58
rect -82 -59 -78 -58
rect -43 -59 -39 -58
rect -2 -59 2 -58
rect 97 -62 101 -50
rect 115 -58 129 -54
rect 153 -57 161 -40
rect 166 -47 170 -32
rect 178 -57 182 -21
rect 209 -22 236 -21
rect 209 -41 213 -22
rect 232 -25 236 -22
rect 256 -28 260 -22
rect 251 -32 260 -28
rect 153 -60 182 -57
rect 187 -46 191 -42
rect 187 -50 197 -46
rect 153 -62 161 -60
rect 187 -62 191 -50
rect 205 -58 219 -54
rect 243 -56 251 -40
rect 256 -47 260 -32
rect 268 -56 272 14
rect 243 -60 272 -56
rect 243 -62 251 -60
rect 137 -66 161 -62
rect 227 -66 251 -62
rect -169 -72 -165 -67
rect -130 -72 -126 -67
rect -90 -72 -86 -67
rect -51 -72 -47 -67
rect -10 -72 -6 -67
rect -173 -76 -153 -72
rect -134 -76 -114 -72
rect -94 -76 -74 -72
rect -55 -76 -35 -72
rect -14 -76 6 -72
rect -187 -92 -163 -88
rect -181 -97 -177 -92
rect -173 -112 -169 -105
rect 122 -99 126 -74
rect 153 -80 161 -66
rect 166 -88 170 -73
rect 161 -92 170 -88
rect 142 -99 146 -95
rect 166 -98 170 -92
rect 122 -103 146 -99
rect 212 -99 216 -74
rect 243 -80 251 -66
rect 256 -88 260 -73
rect 251 -92 260 -88
rect 232 -99 236 -95
rect 256 -98 260 -92
rect 212 -103 236 -99
rect 122 -112 126 -103
rect -195 -116 -188 -112
rect -173 -116 126 -112
rect 212 -112 216 -103
rect 284 -112 288 70
rect 212 -116 288 -112
rect -173 -117 -169 -116
rect -181 -130 -177 -125
rect -185 -134 -165 -130
<< labels >>
rlabel metal1 95 81 95 81 1 gnd
rlabel metal1 164 96 164 96 1 vdd
rlabel metal1 164 46 164 46 1 vdd
rlabel metal1 168 -30 168 -30 1 vdd
rlabel metal1 168 -90 168 -90 1 vdd
rlabel metal1 99 -48 99 -48 1 gnd
rlabel metal1 86 21 86 21 1 vdd
rlabel metal1 86 -21 86 -21 1 gnd
rlabel metal1 63 28 63 28 1 vdd
rlabel metal1 63 -32 63 -32 1 vdd
rlabel metal1 -6 10 -6 10 1 gnd
rlabel metal1 -167 -32 -167 -32 1 vdd
rlabel metal1 -127 -32 -127 -32 1 vdd
rlabel metal1 -128 -74 -128 -74 1 gnd
rlabel metal1 -167 -74 -167 -74 1 gnd
rlabel metal1 -88 -32 -88 -32 1 vdd
rlabel metal1 -88 -74 -88 -74 1 gnd
rlabel metal1 -49 -31 -49 -31 1 vdd
rlabel metal1 -49 -74 -49 -74 1 gnd
rlabel metal1 -8 -31 -8 -31 1 vdd
rlabel metal1 -8 -73 -8 -73 1 gnd
rlabel metal1 -179 -132 -179 -132 1 gnd
rlabel metal1 -180 -90 -180 -90 1 vdd
rlabel metal1 -181 43 -181 43 4 clk
rlabel metal1 185 78 185 78 1 gnd
rlabel metal1 254 40 254 40 1 vdd
rlabel metal1 254 97 254 97 1 vdd
rlabel metal1 189 -48 189 -48 1 gnd
rlabel metal1 258 -90 258 -90 7 vdd
rlabel metal1 258 -30 258 -30 7 vdd
rlabel metal1 258 226 258 226 7 vdd
rlabel metal1 258 166 258 166 7 vdd
rlabel metal1 189 208 189 208 1 gnd
rlabel metal1 254 353 254 353 1 vdd
rlabel metal1 254 296 254 296 1 vdd
rlabel metal1 185 334 185 334 1 gnd
rlabel metal1 -181 299 -181 299 4 clk
rlabel metal1 -180 166 -180 166 1 vdd
rlabel metal1 -179 124 -179 124 1 gnd
rlabel metal1 -8 183 -8 183 1 gnd
rlabel metal1 -8 225 -8 225 1 vdd
rlabel metal1 -49 182 -49 182 1 gnd
rlabel metal1 -49 225 -49 225 1 vdd
rlabel metal1 -88 182 -88 182 1 gnd
rlabel metal1 -88 224 -88 224 1 vdd
rlabel metal1 -167 182 -167 182 1 gnd
rlabel metal1 -128 182 -128 182 1 gnd
rlabel metal1 -127 224 -127 224 1 vdd
rlabel metal1 -167 224 -167 224 1 vdd
rlabel metal1 -6 266 -6 266 1 gnd
rlabel metal1 63 224 63 224 1 vdd
rlabel metal1 63 284 63 284 1 vdd
rlabel metal1 86 235 86 235 1 gnd
rlabel metal1 86 277 86 277 1 vdd
rlabel metal1 99 208 99 208 1 gnd
rlabel metal1 168 166 168 166 1 vdd
rlabel metal1 168 226 168 226 1 vdd
rlabel metal1 164 302 164 302 1 vdd
rlabel metal1 164 352 164 352 1 vdd
rlabel metal1 95 337 95 337 1 gnd
rlabel metal1 258 482 258 482 7 vdd
rlabel metal1 258 422 258 422 7 vdd
rlabel metal1 189 464 189 464 1 gnd
rlabel metal1 254 609 254 609 1 vdd
rlabel metal1 254 552 254 552 1 vdd
rlabel metal1 185 590 185 590 1 gnd
rlabel metal1 -181 555 -181 555 4 clk
rlabel metal1 -180 422 -180 422 1 vdd
rlabel metal1 -179 380 -179 380 1 gnd
rlabel metal1 -8 439 -8 439 1 gnd
rlabel metal1 -8 481 -8 481 1 vdd
rlabel metal1 -49 438 -49 438 1 gnd
rlabel metal1 -49 481 -49 481 1 vdd
rlabel metal1 -88 438 -88 438 1 gnd
rlabel metal1 -88 480 -88 480 1 vdd
rlabel metal1 -167 438 -167 438 1 gnd
rlabel metal1 -128 438 -128 438 1 gnd
rlabel metal1 -127 480 -127 480 1 vdd
rlabel metal1 -167 480 -167 480 1 vdd
rlabel metal1 -6 522 -6 522 1 gnd
rlabel metal1 63 480 63 480 1 vdd
rlabel metal1 63 540 63 540 1 vdd
rlabel metal1 86 491 86 491 1 gnd
rlabel metal1 86 533 86 533 1 vdd
rlabel metal1 99 464 99 464 1 gnd
rlabel metal1 168 422 168 422 1 vdd
rlabel metal1 168 482 168 482 1 vdd
rlabel metal1 164 558 164 558 1 vdd
rlabel metal1 164 608 164 608 1 vdd
rlabel metal1 95 593 95 593 1 gnd
rlabel metal1 258 738 258 738 7 vdd
rlabel metal1 258 678 258 678 7 vdd
rlabel metal1 189 720 189 720 1 gnd
rlabel metal1 254 808 254 808 1 vdd
rlabel metal1 185 846 185 846 1 gnd
rlabel metal1 -181 811 -181 811 4 clk
rlabel metal1 -180 678 -180 678 1 vdd
rlabel metal1 -179 636 -179 636 1 gnd
rlabel metal1 -8 695 -8 695 1 gnd
rlabel metal1 -8 737 -8 737 1 vdd
rlabel metal1 -49 694 -49 694 1 gnd
rlabel metal1 -49 737 -49 737 1 vdd
rlabel metal1 -88 694 -88 694 1 gnd
rlabel metal1 -88 736 -88 736 1 vdd
rlabel metal1 -167 694 -167 694 1 gnd
rlabel metal1 -128 694 -128 694 1 gnd
rlabel metal1 -127 736 -127 736 1 vdd
rlabel metal1 -167 736 -167 736 1 vdd
rlabel metal1 -6 778 -6 778 1 gnd
rlabel metal1 63 736 63 736 1 vdd
rlabel metal1 63 796 63 796 1 vdd
rlabel metal1 86 747 86 747 1 gnd
rlabel metal1 86 789 86 789 1 vdd
rlabel metal1 99 720 99 720 1 gnd
rlabel metal1 168 678 168 678 1 vdd
rlabel metal1 168 738 168 738 1 vdd
rlabel metal1 164 814 164 814 1 vdd
rlabel metal1 164 864 164 864 1 vdd
rlabel metal1 95 849 95 849 1 gnd
rlabel metal1 254 865 254 865 1 vdd
rlabel metal1 95 1105 95 1105 1 gnd
rlabel metal1 164 1120 164 1120 1 vdd
rlabel metal1 164 1070 164 1070 1 vdd
rlabel metal1 168 994 168 994 1 vdd
rlabel metal1 168 934 168 934 1 vdd
rlabel metal1 99 976 99 976 1 gnd
rlabel metal1 86 1045 86 1045 1 vdd
rlabel metal1 86 1003 86 1003 1 gnd
rlabel metal1 63 1052 63 1052 1 vdd
rlabel metal1 63 992 63 992 1 vdd
rlabel metal1 -6 1034 -6 1034 1 gnd
rlabel metal1 -167 992 -167 992 1 vdd
rlabel metal1 -127 992 -127 992 1 vdd
rlabel metal1 -128 950 -128 950 1 gnd
rlabel metal1 -167 950 -167 950 1 gnd
rlabel metal1 -88 992 -88 992 1 vdd
rlabel metal1 -88 950 -88 950 1 gnd
rlabel metal1 -49 993 -49 993 1 vdd
rlabel metal1 -49 950 -49 950 1 gnd
rlabel metal1 -8 993 -8 993 1 vdd
rlabel metal1 -8 951 -8 951 1 gnd
rlabel metal1 -179 892 -179 892 1 gnd
rlabel metal1 -180 934 -180 934 1 vdd
rlabel metal1 -181 1067 -181 1067 4 clk
rlabel metal1 185 1102 185 1102 1 gnd
rlabel metal1 254 1064 254 1064 1 vdd
rlabel metal1 254 1121 254 1121 1 vdd
rlabel metal1 189 976 189 976 1 gnd
rlabel metal1 258 934 258 934 7 vdd
rlabel metal1 258 994 258 994 7 vdd
rlabel metal1 258 1250 258 1250 7 vdd
rlabel metal1 258 1190 258 1190 7 vdd
rlabel metal1 189 1232 189 1232 1 gnd
rlabel metal1 254 1377 254 1377 1 vdd
rlabel metal1 254 1320 254 1320 1 vdd
rlabel metal1 185 1358 185 1358 1 gnd
rlabel metal1 -181 1323 -181 1323 4 clk
rlabel metal1 -180 1190 -180 1190 1 vdd
rlabel metal1 -179 1148 -179 1148 1 gnd
rlabel metal1 -8 1207 -8 1207 1 gnd
rlabel metal1 -8 1249 -8 1249 1 vdd
rlabel metal1 -49 1206 -49 1206 1 gnd
rlabel metal1 -49 1249 -49 1249 1 vdd
rlabel metal1 -88 1206 -88 1206 1 gnd
rlabel metal1 -88 1248 -88 1248 1 vdd
rlabel metal1 -167 1206 -167 1206 1 gnd
rlabel metal1 -128 1206 -128 1206 1 gnd
rlabel metal1 -127 1248 -127 1248 1 vdd
rlabel metal1 -167 1248 -167 1248 1 vdd
rlabel metal1 -6 1290 -6 1290 1 gnd
rlabel metal1 63 1248 63 1248 1 vdd
rlabel metal1 63 1308 63 1308 1 vdd
rlabel metal1 86 1259 86 1259 1 gnd
rlabel metal1 86 1301 86 1301 1 vdd
rlabel metal1 99 1232 99 1232 1 gnd
rlabel metal1 168 1190 168 1190 1 vdd
rlabel metal1 168 1250 168 1250 1 vdd
rlabel metal1 164 1326 164 1326 1 vdd
rlabel metal1 164 1376 164 1376 1 vdd
rlabel metal1 95 1361 95 1361 1 gnd
rlabel metal1 258 1506 258 1506 7 vdd
rlabel metal1 258 1446 258 1446 7 vdd
rlabel metal1 189 1488 189 1488 1 gnd
rlabel metal1 254 1633 254 1633 1 vdd
rlabel metal1 254 1576 254 1576 1 vdd
rlabel metal1 185 1614 185 1614 1 gnd
rlabel metal1 -181 1579 -181 1579 4 clk
rlabel metal1 -180 1446 -180 1446 1 vdd
rlabel metal1 -179 1404 -179 1404 1 gnd
rlabel metal1 -8 1463 -8 1463 1 gnd
rlabel metal1 -8 1505 -8 1505 1 vdd
rlabel metal1 -49 1462 -49 1462 1 gnd
rlabel metal1 -49 1505 -49 1505 1 vdd
rlabel metal1 -88 1462 -88 1462 1 gnd
rlabel metal1 -88 1504 -88 1504 1 vdd
rlabel metal1 -167 1462 -167 1462 1 gnd
rlabel metal1 -128 1462 -128 1462 1 gnd
rlabel metal1 -127 1504 -127 1504 1 vdd
rlabel metal1 -167 1504 -167 1504 1 vdd
rlabel metal1 -6 1546 -6 1546 1 gnd
rlabel metal1 63 1504 63 1504 1 vdd
rlabel metal1 63 1564 63 1564 1 vdd
rlabel metal1 86 1515 86 1515 1 gnd
rlabel metal1 86 1557 86 1557 1 vdd
rlabel metal1 99 1488 99 1488 1 gnd
rlabel metal1 168 1446 168 1446 1 vdd
rlabel metal1 168 1506 168 1506 1 vdd
rlabel metal1 164 1582 164 1582 1 vdd
rlabel metal1 164 1632 164 1632 1 vdd
rlabel metal1 95 1617 95 1617 1 gnd
rlabel metal1 258 1762 258 1762 7 vdd
rlabel metal1 258 1702 258 1702 7 vdd
rlabel metal1 189 1744 189 1744 1 gnd
rlabel metal1 254 1889 254 1889 1 vdd
rlabel metal1 254 1832 254 1832 1 vdd
rlabel metal1 185 1870 185 1870 1 gnd
rlabel metal1 -181 1835 -181 1835 4 clk
rlabel metal1 -180 1702 -180 1702 1 vdd
rlabel metal1 -179 1660 -179 1660 1 gnd
rlabel metal1 -8 1719 -8 1719 1 gnd
rlabel metal1 -8 1761 -8 1761 1 vdd
rlabel metal1 -49 1718 -49 1718 1 gnd
rlabel metal1 -49 1761 -49 1761 1 vdd
rlabel metal1 -88 1718 -88 1718 1 gnd
rlabel metal1 -88 1760 -88 1760 1 vdd
rlabel metal1 -167 1718 -167 1718 1 gnd
rlabel metal1 -128 1718 -128 1718 1 gnd
rlabel metal1 -127 1760 -127 1760 1 vdd
rlabel metal1 -167 1760 -167 1760 1 vdd
rlabel metal1 -6 1802 -6 1802 1 gnd
rlabel metal1 63 1760 63 1760 1 vdd
rlabel metal1 63 1820 63 1820 1 vdd
rlabel metal1 86 1771 86 1771 1 gnd
rlabel metal1 86 1813 86 1813 1 vdd
rlabel metal1 99 1744 99 1744 1 gnd
rlabel metal1 168 1702 168 1702 1 vdd
rlabel metal1 168 1762 168 1762 1 vdd
rlabel metal1 164 1838 164 1838 1 vdd
rlabel metal1 164 1888 164 1888 1 vdd
rlabel metal1 95 1873 95 1873 1 gnd
rlabel metal1 -193 1902 -193 1902 4 a0
rlabel metal1 -193 110 -193 110 3 b3
rlabel metal1 -193 1646 -193 1646 3 b0
rlabel metal1 -193 1390 -193 1390 3 a1
rlabel metal1 -193 1134 -193 1134 3 b1
rlabel metal1 -193 878 -193 878 3 a2
rlabel metal1 -193 622 -193 622 3 b2
rlabel metal1 -193 366 -193 366 3 a3
rlabel metal1 286 1864 286 1864 1 ffa0
rlabel metal1 270 1734 270 1734 1 ffa0_bar
rlabel metal1 286 1608 286 1608 1 ffb0
rlabel metal1 270 1478 270 1478 1 ffb0_bar
rlabel metal1 286 1352 286 1352 1 ffa1
rlabel metal1 270 1222 270 1222 1 ffa1_bar
rlabel metal1 286 1096 286 1096 1 ffb1
rlabel metal1 270 966 270 966 1 ffb1_bar
rlabel metal1 286 840 286 840 1 ffa2
rlabel metal1 270 710 270 710 1 ffa2_bar
rlabel metal1 286 584 286 584 1 ffb2
rlabel metal1 270 454 270 454 1 ffb2_bar
rlabel metal1 286 328 286 328 1 ffa3
rlabel metal1 270 198 270 198 1 ffa3_bar
rlabel metal1 286 72 286 72 1 ffb3
rlabel metal1 270 -58 270 -58 1 ffb3_bar
rlabel metal1 351 476 351 476 1 gnd
rlabel metal1 420 434 420 434 7 vdd
rlabel metal1 420 494 420 494 7 vdd
rlabel metal1 351 381 351 381 1 gnd
rlabel metal1 420 339 420 339 7 vdd
rlabel metal1 420 399 420 399 7 vdd
rlabel metal1 506 449 506 449 7 vdd
rlabel metal1 506 389 506 389 7 vdd
rlabel metal1 437 431 437 431 1 gnd
rlabel metal1 306 268 306 268 1 gnd
rlabel metal1 375 226 375 226 7 vdd
rlabel metal1 375 286 375 286 7 vdd
rlabel metal1 399 240 399 240 1 gnd
rlabel metal1 400 282 400 282 1 vdd
rlabel metal1 351 811 351 811 1 gnd
rlabel metal1 420 769 420 769 7 vdd
rlabel metal1 420 829 420 829 7 vdd
rlabel metal1 351 716 351 716 1 gnd
rlabel metal1 420 674 420 674 7 vdd
rlabel metal1 420 734 420 734 7 vdd
rlabel metal1 506 784 506 784 7 vdd
rlabel metal1 506 724 506 724 7 vdd
rlabel metal1 437 766 437 766 1 gnd
rlabel metal1 306 603 306 603 1 gnd
rlabel metal1 375 561 375 561 7 vdd
rlabel metal1 375 621 375 621 7 vdd
rlabel metal1 399 575 399 575 1 gnd
rlabel metal1 400 617 400 617 1 vdd
rlabel metal1 351 1146 351 1146 1 gnd
rlabel metal1 420 1104 420 1104 7 vdd
rlabel metal1 420 1164 420 1164 7 vdd
rlabel metal1 351 1051 351 1051 1 gnd
rlabel metal1 420 1009 420 1009 7 vdd
rlabel metal1 420 1069 420 1069 7 vdd
rlabel metal1 506 1119 506 1119 7 vdd
rlabel metal1 506 1059 506 1059 7 vdd
rlabel metal1 437 1101 437 1101 1 gnd
rlabel metal1 306 938 306 938 1 gnd
rlabel metal1 375 896 375 896 7 vdd
rlabel metal1 375 956 375 956 7 vdd
rlabel metal1 399 910 399 910 1 gnd
rlabel metal1 400 952 400 952 1 vdd
rlabel metal1 400 1287 400 1287 1 vdd
rlabel metal1 399 1245 399 1245 1 gnd
rlabel metal1 375 1291 375 1291 7 vdd
rlabel metal1 375 1231 375 1231 7 vdd
rlabel metal1 306 1273 306 1273 1 gnd
rlabel metal1 437 1436 437 1436 1 gnd
rlabel metal1 506 1394 506 1394 7 vdd
rlabel metal1 506 1454 506 1454 7 vdd
rlabel metal1 420 1404 420 1404 7 vdd
rlabel metal1 420 1344 420 1344 7 vdd
rlabel metal1 351 1386 351 1386 1 gnd
rlabel metal1 420 1499 420 1499 7 vdd
rlabel metal1 420 1439 420 1439 7 vdd
rlabel metal1 351 1481 351 1481 1 gnd
rlabel metal1 328 1301 328 1301 1 ffa0
rlabel metal1 331 1220 331 1220 1 ffb0
rlabel metal1 328 966 328 966 1 ffa1
rlabel metal1 331 885 331 885 1 ffb1
rlabel metal1 328 631 328 631 1 ffa2
rlabel metal1 331 550 331 550 1 ffb2
rlabel metal1 328 296 328 296 1 ffa3
rlabel metal1 331 215 331 215 1 ffb3
rlabel metal1 504 1426 504 1426 1 p0
rlabel metal1 421 1263 421 1263 1 g0
rlabel metal1 504 1091 504 1091 1 p1
rlabel metal1 421 928 421 928 1 g1
rlabel metal1 504 756 504 756 1 p2
rlabel metal1 421 593 421 593 1 g2
rlabel metal1 504 421 504 421 1 p3
rlabel metal1 421 258 421 258 1 g3
rlabel metal1 544 1038 544 1038 5 vdd
rlabel metal1 582 1038 582 1038 5 vdd
rlabel metal1 620 1038 620 1038 5 vdd
rlabel metal1 658 1038 658 1038 5 vdd
rlabel metal1 528 794 528 794 7 gnd
rlabel metal1 515 1014 515 1014 1 clk_mcc
rlabel metal1 527 845 527 845 1 c_in
rlabel metal1 535 874 535 874 1 p0
rlabel metal1 565 885 565 885 1 g0
rlabel metal1 602 896 602 896 1 p1
rlabel metal1 603 926 603 926 1 g1
rlabel metal1 640 937 640 937 1 p2
rlabel metal1 641 967 641 967 1 g2
rlabel metal1 678 978 678 978 1 p3
rlabel metal1 708 979 708 979 1 g3
rlabel metal1 582 895 582 895 1 c1_bar
rlabel metal1 620 936 620 936 1 c2_bar
rlabel metal1 658 977 658 977 1 c3_bar
rlabel metal1 696 1002 696 1002 1 cout_bar
rlabel metal1 727 997 727 997 1 gnd
rlabel metal1 728 1039 728 1039 1 vdd
rlabel metal1 727 940 727 940 1 gnd
rlabel metal1 728 982 728 982 1 vdd
rlabel metal1 727 883 727 883 1 gnd
rlabel metal1 728 925 728 925 1 vdd
rlabel metal1 727 826 727 826 1 gnd
rlabel metal1 728 868 728 868 1 vdd
rlabel metal1 714 1015 714 1015 1 cout_bar
rlabel metal1 746 1015 746 1015 1 cout
rlabel metal1 714 958 714 958 1 c1_bar
rlabel metal1 746 958 746 958 1 c1
rlabel metal1 714 901 714 901 1 c2_bar
rlabel metal1 746 901 746 901 1 c2
rlabel metal1 714 844 714 844 1 c3_bar
rlabel metal1 746 844 746 844 1 c3
rlabel metal1 897 1061 897 1061 1 gnd
rlabel metal1 966 1019 966 1019 7 vdd
rlabel metal1 966 1079 966 1079 7 vdd
rlabel metal1 880 1029 880 1029 7 vdd
rlabel metal1 880 969 880 969 7 vdd
rlabel metal1 811 1011 811 1011 1 gnd
rlabel metal1 880 1124 880 1124 7 vdd
rlabel metal1 880 1064 880 1064 7 vdd
rlabel metal1 811 1106 811 1106 1 gnd
rlabel metal1 897 828 897 828 1 gnd
rlabel metal1 966 786 966 786 7 vdd
rlabel metal1 966 846 966 846 7 vdd
rlabel metal1 880 796 880 796 7 vdd
rlabel metal1 880 736 880 736 7 vdd
rlabel metal1 811 778 811 778 1 gnd
rlabel metal1 880 891 880 891 7 vdd
rlabel metal1 880 831 880 831 7 vdd
rlabel metal1 811 873 811 873 1 gnd
rlabel metal1 811 1339 811 1339 1 gnd
rlabel metal1 880 1297 880 1297 7 vdd
rlabel metal1 880 1357 880 1357 7 vdd
rlabel metal1 811 1244 811 1244 1 gnd
rlabel metal1 880 1202 880 1202 7 vdd
rlabel metal1 880 1262 880 1262 7 vdd
rlabel metal1 966 1312 966 1312 7 vdd
rlabel metal1 966 1252 966 1252 7 vdd
rlabel metal1 897 1294 897 1294 1 gnd
rlabel metal1 897 595 897 595 1 gnd
rlabel metal1 966 553 966 553 7 vdd
rlabel metal1 966 613 966 613 7 vdd
rlabel metal1 880 563 880 563 7 vdd
rlabel metal1 880 503 880 503 7 vdd
rlabel metal1 811 545 811 545 1 gnd
rlabel metal1 880 658 880 658 7 vdd
rlabel metal1 880 598 880 598 7 vdd
rlabel metal1 811 640 811 640 1 gnd
rlabel metal1 782 474 782 474 1 gnd
rlabel metal1 783 516 783 516 1 vdd
rlabel metal1 360 1426 360 1426 3 vdd
rlabel metal1 318 1427 318 1427 3 gnd
rlabel metal1 318 1092 318 1092 3 gnd
rlabel metal1 360 1091 360 1091 3 vdd
rlabel metal1 360 756 360 756 3 vdd
rlabel metal1 318 757 318 757 3 gnd
rlabel metal1 360 421 360 421 3 vdd
rlabel metal1 318 422 318 422 3 gnd
rlabel metal1 778 1285 778 1285 3 gnd
rlabel metal1 820 1284 820 1284 3 vdd
rlabel metal1 778 1052 778 1052 3 gnd
rlabel metal1 820 1051 820 1051 3 vdd
rlabel metal1 778 819 778 819 3 gnd
rlabel metal1 820 818 820 818 3 vdd
rlabel metal1 778 586 778 586 3 gnd
rlabel metal1 820 585 820 585 3 vdd
rlabel metal1 322 1491 322 1491 1 gnd
rlabel metal1 323 1533 323 1533 1 vdd
rlabel metal1 322 1156 322 1156 1 gnd
rlabel metal1 323 1198 323 1198 1 vdd
rlabel metal1 323 863 323 863 1 vdd
rlabel metal1 322 821 322 821 1 gnd
rlabel metal1 323 528 323 528 1 vdd
rlabel metal1 322 486 322 486 1 gnd
rlabel metal1 783 1391 783 1391 1 vdd
rlabel metal1 782 1349 782 1349 1 gnd
rlabel metal1 782 1116 782 1116 1 gnd
rlabel metal1 783 1158 783 1158 1 vdd
rlabel metal1 782 883 782 883 1 gnd
rlabel metal1 783 925 783 925 1 vdd
rlabel metal1 782 650 782 650 1 gnd
rlabel metal1 783 692 783 692 1 vdd
rlabel metal1 306 1509 306 1509 1 ffa0
rlabel metal1 336 1442 336 1442 1 ffb0
rlabel metal1 306 1174 306 1174 1 ffa1
rlabel metal1 336 1107 336 1107 1 ffb1
rlabel metal1 306 839 306 839 1 ffa2
rlabel metal1 336 772 336 772 1 ffb2
rlabel metal1 306 504 306 504 1 ffa3
rlabel metal1 336 437 336 437 1 ffb3
rlabel metal1 766 1367 766 1367 1 p0
rlabel metal1 796 1300 796 1300 1 cin
rlabel metal1 766 1134 766 1134 1 p1
rlabel metal1 796 1067 796 1067 1 c1
rlabel metal1 766 901 766 901 1 p2
rlabel metal1 796 834 796 834 1 c2
rlabel metal1 766 668 766 668 1 p3
rlabel metal1 796 601 796 601 1 c3
rlabel metal1 966 585 966 585 1 s3
rlabel metal1 966 818 966 818 1 s2
rlabel metal1 966 1051 966 1051 1 s1
rlabel metal1 966 1284 966 1284 1 s0
rlabel metal1 1277 494 1277 494 1 gnd
rlabel metal1 1346 509 1346 509 1 vdd
rlabel metal1 1346 459 1346 459 1 vdd
rlabel metal1 1350 383 1350 383 1 vdd
rlabel metal1 1350 323 1350 323 1 vdd
rlabel metal1 1281 365 1281 365 1 gnd
rlabel metal1 1268 434 1268 434 1 vdd
rlabel metal1 1268 392 1268 392 1 gnd
rlabel metal1 1245 441 1245 441 1 vdd
rlabel metal1 1245 381 1245 381 1 vdd
rlabel metal1 1176 423 1176 423 1 gnd
rlabel metal1 1015 381 1015 381 1 vdd
rlabel metal1 1055 381 1055 381 1 vdd
rlabel metal1 1054 339 1054 339 1 gnd
rlabel metal1 1015 339 1015 339 1 gnd
rlabel metal1 1094 381 1094 381 1 vdd
rlabel metal1 1094 339 1094 339 1 gnd
rlabel metal1 1133 382 1133 382 1 vdd
rlabel metal1 1133 339 1133 339 1 gnd
rlabel metal1 1174 382 1174 382 1 vdd
rlabel metal1 1174 340 1174 340 1 gnd
rlabel metal1 1003 281 1003 281 1 gnd
rlabel metal1 1002 323 1002 323 1 vdd
rlabel metal1 1001 456 1001 456 4 clk
rlabel metal1 1367 491 1367 491 1 gnd
rlabel metal1 1436 453 1436 453 1 vdd
rlabel metal1 1436 510 1436 510 1 vdd
rlabel metal1 1371 365 1371 365 1 gnd
rlabel metal1 1440 323 1440 323 7 vdd
rlabel metal1 1440 383 1440 383 7 vdd
rlabel metal1 1440 639 1440 639 7 vdd
rlabel metal1 1440 579 1440 579 7 vdd
rlabel metal1 1371 621 1371 621 1 gnd
rlabel metal1 1436 766 1436 766 1 vdd
rlabel metal1 1436 709 1436 709 1 vdd
rlabel metal1 1367 747 1367 747 1 gnd
rlabel metal1 1001 712 1001 712 4 clk
rlabel metal1 1002 579 1002 579 1 vdd
rlabel metal1 1003 537 1003 537 1 gnd
rlabel metal1 1174 596 1174 596 1 gnd
rlabel metal1 1174 638 1174 638 1 vdd
rlabel metal1 1133 595 1133 595 1 gnd
rlabel metal1 1133 638 1133 638 1 vdd
rlabel metal1 1094 595 1094 595 1 gnd
rlabel metal1 1094 637 1094 637 1 vdd
rlabel metal1 1015 595 1015 595 1 gnd
rlabel metal1 1054 595 1054 595 1 gnd
rlabel metal1 1055 637 1055 637 1 vdd
rlabel metal1 1015 637 1015 637 1 vdd
rlabel metal1 1176 679 1176 679 1 gnd
rlabel metal1 1245 637 1245 637 1 vdd
rlabel metal1 1245 697 1245 697 1 vdd
rlabel metal1 1268 648 1268 648 1 gnd
rlabel metal1 1268 690 1268 690 1 vdd
rlabel metal1 1281 621 1281 621 1 gnd
rlabel metal1 1350 579 1350 579 1 vdd
rlabel metal1 1350 639 1350 639 1 vdd
rlabel metal1 1346 715 1346 715 1 vdd
rlabel metal1 1346 765 1346 765 1 vdd
rlabel metal1 1277 750 1277 750 1 gnd
rlabel metal1 1440 895 1440 895 7 vdd
rlabel metal1 1440 835 1440 835 7 vdd
rlabel metal1 1371 877 1371 877 1 gnd
rlabel metal1 1436 1022 1436 1022 1 vdd
rlabel metal1 1436 965 1436 965 1 vdd
rlabel metal1 1367 1003 1367 1003 1 gnd
rlabel metal1 1001 968 1001 968 4 clk
rlabel metal1 1002 835 1002 835 1 vdd
rlabel metal1 1003 793 1003 793 1 gnd
rlabel metal1 1174 852 1174 852 1 gnd
rlabel metal1 1174 894 1174 894 1 vdd
rlabel metal1 1133 851 1133 851 1 gnd
rlabel metal1 1133 894 1133 894 1 vdd
rlabel metal1 1094 851 1094 851 1 gnd
rlabel metal1 1094 893 1094 893 1 vdd
rlabel metal1 1015 851 1015 851 1 gnd
rlabel metal1 1054 851 1054 851 1 gnd
rlabel metal1 1055 893 1055 893 1 vdd
rlabel metal1 1015 893 1015 893 1 vdd
rlabel metal1 1176 935 1176 935 1 gnd
rlabel metal1 1245 893 1245 893 1 vdd
rlabel metal1 1245 953 1245 953 1 vdd
rlabel metal1 1268 904 1268 904 1 gnd
rlabel metal1 1268 946 1268 946 1 vdd
rlabel metal1 1281 877 1281 877 1 gnd
rlabel metal1 1350 835 1350 835 1 vdd
rlabel metal1 1350 895 1350 895 1 vdd
rlabel metal1 1346 971 1346 971 1 vdd
rlabel metal1 1346 1021 1346 1021 1 vdd
rlabel metal1 1277 1006 1277 1006 1 gnd
rlabel metal1 1440 1151 1440 1151 7 vdd
rlabel metal1 1440 1091 1440 1091 7 vdd
rlabel metal1 1371 1133 1371 1133 1 gnd
rlabel metal1 1436 1221 1436 1221 1 vdd
rlabel metal1 1367 1259 1367 1259 1 gnd
rlabel metal1 1001 1224 1001 1224 4 clk
rlabel metal1 1002 1091 1002 1091 1 vdd
rlabel metal1 1003 1049 1003 1049 1 gnd
rlabel metal1 1174 1108 1174 1108 1 gnd
rlabel metal1 1174 1150 1174 1150 1 vdd
rlabel metal1 1133 1107 1133 1107 1 gnd
rlabel metal1 1133 1150 1133 1150 1 vdd
rlabel metal1 1094 1107 1094 1107 1 gnd
rlabel metal1 1094 1149 1094 1149 1 vdd
rlabel metal1 1015 1107 1015 1107 1 gnd
rlabel metal1 1054 1107 1054 1107 1 gnd
rlabel metal1 1055 1149 1055 1149 1 vdd
rlabel metal1 1015 1149 1015 1149 1 vdd
rlabel metal1 1176 1191 1176 1191 1 gnd
rlabel metal1 1245 1149 1245 1149 1 vdd
rlabel metal1 1245 1209 1245 1209 1 vdd
rlabel metal1 1268 1160 1268 1160 1 gnd
rlabel metal1 1268 1202 1268 1202 1 vdd
rlabel metal1 1281 1133 1281 1133 1 gnd
rlabel metal1 1350 1091 1350 1091 1 vdd
rlabel metal1 1350 1151 1350 1151 1 vdd
rlabel metal1 1346 1227 1346 1227 1 vdd
rlabel metal1 1346 1277 1346 1277 1 vdd
rlabel metal1 1277 1262 1277 1262 1 gnd
rlabel metal1 1436 1278 1436 1278 1 vdd
rlabel metal1 1277 1518 1277 1518 1 gnd
rlabel metal1 1346 1533 1346 1533 1 vdd
rlabel metal1 1346 1483 1346 1483 1 vdd
rlabel metal1 1350 1407 1350 1407 1 vdd
rlabel metal1 1350 1347 1350 1347 1 vdd
rlabel metal1 1281 1389 1281 1389 1 gnd
rlabel metal1 1268 1458 1268 1458 1 vdd
rlabel metal1 1268 1416 1268 1416 1 gnd
rlabel metal1 1245 1465 1245 1465 1 vdd
rlabel metal1 1245 1405 1245 1405 1 vdd
rlabel metal1 1176 1447 1176 1447 1 gnd
rlabel metal1 1015 1405 1015 1405 1 vdd
rlabel metal1 1055 1405 1055 1405 1 vdd
rlabel metal1 1054 1363 1054 1363 1 gnd
rlabel metal1 1015 1363 1015 1363 1 gnd
rlabel metal1 1094 1405 1094 1405 1 vdd
rlabel metal1 1094 1363 1094 1363 1 gnd
rlabel metal1 1133 1406 1133 1406 1 vdd
rlabel metal1 1133 1363 1133 1363 1 gnd
rlabel metal1 1174 1406 1174 1406 1 vdd
rlabel metal1 1174 1364 1174 1364 1 gnd
rlabel metal1 1003 1305 1003 1305 1 gnd
rlabel metal1 1002 1347 1002 1347 1 vdd
rlabel metal1 1001 1480 1001 1480 4 clk
rlabel metal1 1367 1515 1367 1515 1 gnd
rlabel metal1 1436 1477 1436 1477 1 vdd
rlabel metal1 1436 1534 1436 1534 1 vdd
rlabel metal1 1371 1389 1371 1389 1 gnd
rlabel metal1 1440 1347 1440 1347 7 vdd
rlabel metal1 1440 1407 1440 1407 7 vdd
rlabel metal1 989 1547 989 1547 1 cout
rlabel metal1 989 1291 989 1291 1 s0
rlabel metal1 989 1035 989 1035 1 s1
rlabel metal1 989 779 989 779 1 s2
rlabel metal1 989 523 989 523 1 s3
rlabel metal1 1468 1509 1468 1509 7 ffcout
rlabel metal1 1452 1379 1452 1379 1 ffcout_bar
rlabel metal1 1468 1253 1468 1253 7 ffs0
rlabel metal1 1452 1123 1452 1123 1 ffs0_bar
rlabel metal1 1468 997 1468 997 7 ffs1
rlabel metal1 1452 867 1452 867 1 ffs1_bar
rlabel metal1 1468 741 1468 741 7 ffs2
rlabel metal1 1452 611 1452 611 1 ffs2_bar
rlabel metal1 1468 485 1468 485 7 ffs3
rlabel metal1 1452 355 1452 355 1 ffs3_bar
<< end >>
