magic
tech scmos
timestamp 1618921300
<< nwell >>
rect 143 83 169 109
rect 233 83 259 109
rect 42 11 68 37
rect 143 31 169 57
rect 233 31 259 57
rect 77 0 103 26
rect -176 -53 -150 -27
rect -137 -53 -111 -27
rect -97 -53 -71 -27
rect -58 -53 -32 -27
rect -17 -53 9 -27
rect 42 -41 68 -15
rect 147 -47 173 -21
rect 237 -47 263 -21
rect -188 -111 -162 -85
rect 147 -99 173 -73
rect 237 -99 263 -73
<< ntransistor >>
rect 103 77 111 79
rect 193 77 201 79
rect 125 69 133 71
rect 215 69 223 71
rect 2 5 10 7
rect 24 -3 32 -1
rect 89 -14 91 -6
rect 107 -53 115 -51
rect 197 -53 205 -51
rect -164 -67 -162 -59
rect -125 -67 -123 -59
rect -85 -67 -83 -59
rect -46 -67 -44 -59
rect -5 -67 -3 -59
rect 129 -61 137 -59
rect 219 -61 227 -59
rect -176 -125 -174 -117
<< ptransistor >>
rect 149 95 157 97
rect 239 95 247 97
rect 149 43 157 45
rect 239 43 247 45
rect 48 23 56 25
rect 89 6 91 14
rect 48 -29 56 -27
rect 153 -35 161 -33
rect 243 -35 251 -33
rect -164 -47 -162 -39
rect -125 -47 -123 -39
rect -85 -47 -83 -39
rect -46 -47 -44 -39
rect -5 -47 -3 -39
rect 153 -87 161 -85
rect 243 -87 251 -85
rect -176 -105 -174 -97
<< ndiffusion >>
rect 103 79 111 80
rect 193 79 201 80
rect 103 76 111 77
rect 193 76 201 77
rect 125 71 133 72
rect 215 71 223 72
rect 125 68 133 69
rect 215 68 223 69
rect 2 7 10 8
rect 2 4 10 5
rect 24 -1 32 0
rect 24 -4 32 -3
rect 88 -14 89 -6
rect 91 -14 92 -6
rect 107 -51 115 -50
rect 197 -51 205 -50
rect 107 -54 115 -53
rect 197 -54 205 -53
rect 129 -59 137 -58
rect 219 -59 227 -58
rect -165 -67 -164 -59
rect -162 -67 -161 -59
rect -126 -67 -125 -59
rect -123 -67 -122 -59
rect -86 -67 -85 -59
rect -83 -67 -82 -59
rect -47 -67 -46 -59
rect -44 -67 -43 -59
rect -6 -67 -5 -59
rect -3 -67 -2 -59
rect 129 -62 137 -61
rect 219 -62 227 -61
rect -177 -125 -176 -117
rect -174 -125 -173 -117
<< pdiffusion >>
rect 149 97 157 98
rect 239 97 247 98
rect 149 94 157 95
rect 239 94 247 95
rect 149 45 157 46
rect 239 45 247 46
rect 149 42 157 43
rect 239 42 247 43
rect 48 25 56 26
rect 48 22 56 23
rect 88 6 89 14
rect 91 6 92 14
rect 48 -27 56 -26
rect 48 -30 56 -29
rect 153 -33 161 -32
rect 243 -33 251 -32
rect 153 -36 161 -35
rect -165 -47 -164 -39
rect -162 -47 -161 -39
rect -126 -47 -125 -39
rect -123 -47 -122 -39
rect -86 -47 -85 -39
rect -83 -47 -82 -39
rect -47 -47 -46 -39
rect -44 -47 -43 -39
rect -6 -47 -5 -39
rect -3 -47 -2 -39
rect 243 -36 251 -35
rect 153 -85 161 -84
rect 243 -85 251 -84
rect 153 -88 161 -87
rect 243 -88 251 -87
rect -177 -105 -176 -97
rect -174 -105 -173 -97
<< ndcontact >>
rect 103 80 111 84
rect 193 80 201 84
rect 103 72 111 76
rect 125 72 133 76
rect 193 72 201 76
rect 215 72 223 76
rect 125 64 133 68
rect 215 64 223 68
rect 2 8 10 12
rect 2 0 10 4
rect 24 0 32 4
rect 24 -8 32 -4
rect 84 -14 88 -6
rect 92 -14 96 -6
rect 107 -50 115 -46
rect 197 -50 205 -46
rect 107 -58 115 -54
rect 129 -58 137 -54
rect 197 -58 205 -54
rect 219 -58 227 -54
rect -169 -67 -165 -59
rect -161 -67 -157 -59
rect -130 -67 -126 -59
rect -122 -67 -118 -59
rect -90 -67 -86 -59
rect -82 -67 -78 -59
rect -51 -67 -47 -59
rect -43 -67 -39 -59
rect -10 -67 -6 -59
rect -2 -67 2 -59
rect 129 -66 137 -62
rect 219 -66 227 -62
rect -181 -125 -177 -117
rect -173 -125 -169 -117
<< pdcontact >>
rect 149 98 157 102
rect 239 98 247 102
rect 149 90 157 94
rect 239 90 247 94
rect 149 46 157 50
rect 239 46 247 50
rect 149 38 157 42
rect 239 38 247 42
rect 48 26 56 30
rect 48 18 56 22
rect 84 6 88 14
rect 92 6 96 14
rect 48 -26 56 -22
rect 48 -34 56 -30
rect 153 -32 161 -28
rect 243 -32 251 -28
rect -169 -47 -165 -39
rect -161 -47 -157 -39
rect -130 -47 -126 -39
rect -122 -47 -118 -39
rect -90 -47 -86 -39
rect -82 -47 -78 -39
rect -51 -47 -47 -39
rect -43 -47 -39 -39
rect -10 -47 -6 -39
rect -2 -47 2 -39
rect 153 -40 161 -36
rect 243 -40 251 -36
rect 153 -84 161 -80
rect 243 -84 251 -80
rect 153 -92 161 -88
rect 243 -92 251 -88
rect -181 -105 -177 -97
rect -173 -105 -169 -97
<< polysilicon >>
rect 139 97 141 101
rect 229 97 231 101
rect 136 95 149 97
rect 157 95 160 97
rect 226 95 239 97
rect 247 95 250 97
rect 116 79 118 85
rect 206 79 208 85
rect 100 77 103 79
rect 111 77 121 79
rect 190 77 193 79
rect 201 77 211 79
rect 115 69 125 71
rect 133 69 136 71
rect 205 69 215 71
rect 223 69 226 71
rect 119 60 121 69
rect 209 60 211 69
rect 136 43 149 45
rect 157 43 160 45
rect 226 43 239 45
rect 247 43 250 45
rect 139 39 141 43
rect 229 39 231 43
rect 38 25 40 29
rect 35 23 48 25
rect 56 23 59 25
rect 89 14 91 17
rect 15 7 17 13
rect -1 5 2 7
rect 10 5 20 7
rect 14 -3 24 -1
rect 32 -3 35 -1
rect 18 -12 20 -3
rect 89 -2 91 6
rect 81 -4 91 -2
rect 89 -6 91 -4
rect 89 -17 91 -14
rect 35 -29 48 -27
rect 56 -29 59 -27
rect 38 -33 40 -29
rect -164 -39 -162 -36
rect -125 -39 -123 -36
rect -85 -39 -83 -36
rect -46 -39 -44 -36
rect -5 -39 -3 -36
rect 143 -33 145 -29
rect 233 -33 235 -29
rect 140 -35 153 -33
rect 161 -35 164 -33
rect 230 -35 243 -33
rect 251 -35 254 -33
rect -164 -55 -162 -47
rect -172 -57 -162 -55
rect -164 -59 -162 -57
rect -125 -55 -123 -47
rect -133 -57 -123 -55
rect -125 -59 -123 -57
rect -85 -55 -83 -47
rect -93 -57 -83 -55
rect -85 -59 -83 -57
rect -46 -55 -44 -47
rect -54 -57 -44 -55
rect -46 -59 -44 -57
rect -5 -55 -3 -47
rect 120 -51 122 -45
rect 210 -51 212 -45
rect 104 -53 107 -51
rect 115 -53 125 -51
rect 194 -53 197 -51
rect 205 -53 215 -51
rect -13 -57 -3 -55
rect -5 -59 -3 -57
rect 119 -61 129 -59
rect 137 -61 140 -59
rect 209 -61 219 -59
rect 227 -61 230 -59
rect -164 -70 -162 -67
rect -125 -70 -123 -67
rect -85 -70 -83 -67
rect -46 -70 -44 -67
rect -5 -70 -3 -67
rect 123 -70 125 -61
rect 213 -70 215 -61
rect 140 -87 153 -85
rect 161 -87 164 -85
rect 230 -87 243 -85
rect 251 -87 254 -85
rect 143 -91 145 -87
rect -176 -97 -174 -94
rect 233 -91 235 -87
rect -176 -113 -174 -105
rect -184 -115 -174 -113
rect -176 -117 -174 -115
rect -176 -128 -174 -125
<< polycontact >>
rect 138 101 142 105
rect 228 101 232 105
rect 115 85 119 89
rect 205 85 209 89
rect 118 56 122 60
rect 208 56 212 60
rect 138 35 142 39
rect 228 35 232 39
rect 37 29 41 33
rect 14 13 18 17
rect 77 -5 81 -1
rect 17 -16 21 -12
rect 142 -29 146 -25
rect 37 -37 41 -33
rect 232 -29 236 -25
rect 119 -45 123 -41
rect 209 -45 213 -41
rect -176 -58 -172 -54
rect -137 -58 -133 -54
rect -97 -58 -93 -54
rect -58 -58 -54 -54
rect -17 -58 -13 -54
rect 122 -74 126 -70
rect 212 -74 216 -70
rect 142 -95 146 -91
rect 232 -95 236 -91
rect -188 -116 -184 -112
<< metal1 >>
rect -195 108 142 112
rect 174 108 232 112
rect -195 -112 -191 108
rect 115 89 119 108
rect 138 105 142 108
rect 162 102 166 108
rect 157 98 166 102
rect 93 84 97 88
rect 93 80 103 84
rect 93 68 97 80
rect 111 72 125 76
rect 149 74 157 90
rect 162 83 166 98
rect 174 74 178 108
rect 205 89 209 108
rect 228 105 232 108
rect 252 102 256 108
rect 247 98 256 102
rect 149 70 178 74
rect 183 84 187 88
rect 183 80 193 84
rect 149 68 157 70
rect 183 68 187 80
rect 201 72 215 76
rect 239 74 247 90
rect 252 83 256 98
rect 239 70 288 74
rect 239 68 247 70
rect 133 64 157 68
rect 223 64 247 68
rect -183 41 18 45
rect -183 -54 -179 41
rect 14 40 18 41
rect 14 36 41 40
rect 14 17 18 36
rect 37 33 41 36
rect 61 30 65 36
rect 56 26 65 30
rect -8 12 -4 16
rect -8 8 2 12
rect -8 -4 -4 8
rect 10 0 24 4
rect 48 -1 56 18
rect 61 11 65 26
rect 118 31 122 56
rect 149 50 157 64
rect 162 42 166 57
rect 157 38 166 42
rect 138 31 142 35
rect 162 32 166 38
rect 118 27 142 31
rect 208 31 212 56
rect 239 50 247 64
rect 252 42 256 57
rect 247 38 256 42
rect 228 31 232 35
rect 252 32 256 38
rect 208 27 232 31
rect 78 19 102 23
rect 84 14 88 19
rect 92 -1 96 6
rect 118 -1 122 27
rect 208 18 212 27
rect 208 14 272 18
rect 48 -4 77 -1
rect 32 -5 77 -4
rect 92 -5 123 -1
rect 32 -8 56 -5
rect 92 -6 96 -5
rect -175 -34 -151 -30
rect -136 -34 -112 -30
rect -96 -34 -72 -30
rect -57 -34 -33 -30
rect -16 -34 8 -30
rect -169 -39 -165 -34
rect -130 -39 -126 -34
rect -90 -39 -86 -34
rect -51 -39 -47 -34
rect -10 -39 -6 -34
rect -161 -54 -157 -47
rect -122 -54 -118 -47
rect -82 -54 -78 -47
rect -43 -54 -39 -47
rect -2 -54 2 -47
rect 17 -41 21 -16
rect 48 -22 56 -8
rect 61 -30 65 -15
rect 84 -19 88 -14
rect 119 -18 123 -5
rect 80 -23 100 -19
rect 119 -22 146 -18
rect 178 -21 236 -18
rect 56 -34 65 -30
rect 37 -41 41 -37
rect 61 -40 65 -34
rect 17 -45 41 -41
rect 119 -41 123 -22
rect 142 -25 146 -22
rect 166 -28 170 -22
rect 161 -32 170 -28
rect 17 -54 21 -45
rect -183 -58 -176 -54
rect -161 -58 -137 -54
rect -122 -58 -97 -54
rect -82 -58 -58 -54
rect -43 -58 -17 -54
rect -2 -58 21 -54
rect 97 -46 101 -42
rect 97 -50 107 -46
rect -161 -59 -157 -58
rect -122 -59 -118 -58
rect -82 -59 -78 -58
rect -43 -59 -39 -58
rect -2 -59 2 -58
rect 97 -62 101 -50
rect 115 -58 129 -54
rect 153 -57 161 -40
rect 166 -47 170 -32
rect 178 -57 182 -21
rect 209 -22 236 -21
rect 209 -41 213 -22
rect 232 -25 236 -22
rect 256 -28 260 -22
rect 251 -32 260 -28
rect 153 -60 182 -57
rect 187 -46 191 -42
rect 187 -50 197 -46
rect 153 -62 161 -60
rect 187 -62 191 -50
rect 205 -58 219 -54
rect 243 -56 251 -40
rect 256 -47 260 -32
rect 268 -56 272 14
rect 243 -60 272 -56
rect 243 -62 251 -60
rect 137 -66 161 -62
rect 227 -66 251 -62
rect -169 -72 -165 -67
rect -130 -72 -126 -67
rect -90 -72 -86 -67
rect -51 -72 -47 -67
rect -10 -72 -6 -67
rect -173 -76 -153 -72
rect -134 -76 -114 -72
rect -94 -76 -74 -72
rect -55 -76 -35 -72
rect -14 -76 6 -72
rect -187 -92 -163 -88
rect -181 -97 -177 -92
rect -173 -112 -169 -105
rect 122 -99 126 -74
rect 153 -80 161 -66
rect 166 -88 170 -73
rect 161 -92 170 -88
rect 142 -99 146 -95
rect 166 -98 170 -92
rect 122 -103 146 -99
rect 212 -99 216 -74
rect 243 -80 251 -66
rect 256 -88 260 -73
rect 251 -92 260 -88
rect 232 -99 236 -95
rect 256 -98 260 -92
rect 212 -103 236 -99
rect 122 -112 126 -103
rect -195 -116 -188 -112
rect -173 -116 126 -112
rect 212 -112 216 -103
rect 284 -112 288 70
rect 212 -116 288 -112
rect -173 -117 -169 -116
rect -181 -130 -177 -125
rect -185 -134 -165 -130
<< labels >>
rlabel metal1 95 81 95 81 1 gnd
rlabel metal1 164 96 164 96 1 vdd
rlabel metal1 164 46 164 46 1 vdd
rlabel metal1 168 -30 168 -30 1 vdd
rlabel metal1 168 -90 168 -90 1 vdd
rlabel metal1 99 -48 99 -48 1 gnd
rlabel metal1 86 21 86 21 1 vdd
rlabel metal1 86 -21 86 -21 1 gnd
rlabel metal1 63 28 63 28 1 vdd
rlabel metal1 63 -32 63 -32 1 vdd
rlabel metal1 -6 10 -6 10 1 gnd
rlabel metal1 -167 -32 -167 -32 1 vdd
rlabel metal1 -127 -32 -127 -32 1 vdd
rlabel metal1 -128 -74 -128 -74 1 gnd
rlabel metal1 -167 -74 -167 -74 1 gnd
rlabel metal1 -88 -32 -88 -32 1 vdd
rlabel metal1 -88 -74 -88 -74 1 gnd
rlabel metal1 -49 -31 -49 -31 1 vdd
rlabel metal1 -49 -74 -49 -74 1 gnd
rlabel metal1 -8 -31 -8 -31 1 vdd
rlabel metal1 -8 -73 -8 -73 1 gnd
rlabel metal1 -179 -132 -179 -132 1 gnd
rlabel metal1 -180 -90 -180 -90 1 vdd
rlabel metal1 -181 43 -181 43 4 clk
rlabel metal1 -193 110 -193 110 4 d
rlabel metal1 185 78 185 78 1 gnd
rlabel metal1 254 40 254 40 1 vdd
rlabel metal1 254 97 254 97 1 vdd
rlabel metal1 189 -48 189 -48 1 gnd
rlabel metal1 258 -90 258 -90 7 vdd
rlabel metal1 258 -30 258 -30 7 vdd
rlabel metal1 270 -58 270 -58 1 q_bar
rlabel metal1 286 72 286 72 7 q
<< end >>
