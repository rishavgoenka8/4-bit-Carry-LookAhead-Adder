magic
tech scmos
timestamp 1618792186
<< nwell >>
rect 0 0 26 26
<< ntransistor >>
rect 12 -14 14 -6
<< ptransistor >>
rect 12 6 14 14
<< ndiffusion >>
rect 11 -14 12 -6
rect 14 -14 15 -6
<< pdiffusion >>
rect 11 6 12 14
rect 14 6 15 14
<< ndcontact >>
rect 7 -14 11 -6
rect 15 -14 19 -6
<< pdcontact >>
rect 7 6 11 14
rect 15 6 19 14
<< polysilicon >>
rect 12 14 14 17
rect 12 -2 14 6
rect 4 -4 14 -2
rect 12 -6 14 -4
rect 12 -17 14 -14
<< polycontact >>
rect 0 -5 4 -1
<< metal1 >>
rect 1 19 25 22
rect 7 14 11 19
rect 15 -1 19 6
rect -2 -5 0 -1
rect 15 -5 23 -1
rect 15 -6 19 -5
rect 7 -19 11 -14
rect 3 -23 23 -19
<< labels >>
rlabel metal1 6 21 6 21 5 vdd
rlabel metal1 -1 -3 -1 -3 3 in
rlabel metal1 21 -3 21 -3 7 out
rlabel metal1 8 -21 8 -21 1 gnd
<< end >>
