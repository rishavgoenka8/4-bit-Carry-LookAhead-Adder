magic
tech scmos
timestamp 1619593377
<< nwell >>
rect -123 1952 -97 1978
rect -33 1952 -7 1978
rect 143 1951 169 1977
rect 233 1951 259 1977
rect -123 1900 -97 1926
rect -33 1900 -7 1926
rect 143 1899 169 1925
rect 233 1899 259 1925
rect -189 1869 -163 1895
rect -119 1822 -93 1848
rect -29 1822 -3 1848
rect 147 1821 173 1847
rect 237 1821 263 1847
rect -178 1773 -152 1799
rect -119 1770 -93 1796
rect -29 1770 -3 1796
rect 88 1772 114 1798
rect 147 1769 173 1795
rect 237 1769 263 1795
rect -178 1721 -152 1747
rect 88 1720 114 1746
rect -123 1680 -97 1706
rect -33 1680 -7 1706
rect 143 1679 169 1705
rect 233 1679 259 1705
rect -123 1628 -97 1654
rect -33 1628 -7 1654
rect 143 1627 169 1653
rect 233 1627 259 1653
rect -189 1597 -163 1623
rect 1100 1580 1126 1606
rect 1190 1580 1216 1606
rect 1366 1579 1392 1605
rect 1456 1579 1482 1605
rect -119 1550 -93 1576
rect -29 1550 -3 1576
rect 147 1549 173 1575
rect 237 1549 263 1575
rect -178 1501 -152 1527
rect -119 1498 -93 1524
rect -29 1498 -3 1524
rect 88 1500 114 1526
rect 147 1497 173 1523
rect 237 1497 263 1523
rect 313 1512 339 1538
rect 1100 1528 1126 1554
rect 1190 1528 1216 1554
rect 1366 1527 1392 1553
rect 1456 1527 1482 1553
rect 399 1482 425 1508
rect 1034 1497 1060 1523
rect -178 1449 -152 1475
rect 88 1448 114 1474
rect -123 1408 -97 1434
rect -33 1408 -7 1434
rect 143 1407 169 1433
rect 233 1407 259 1433
rect 339 1410 365 1436
rect 399 1430 425 1456
rect 485 1437 511 1463
rect 1104 1450 1130 1476
rect 1194 1450 1220 1476
rect 1370 1449 1396 1475
rect 1460 1449 1486 1475
rect 399 1387 425 1413
rect 485 1385 511 1411
rect 1045 1401 1071 1427
rect 1104 1398 1130 1424
rect 1194 1398 1220 1424
rect 1311 1400 1337 1426
rect 1370 1397 1396 1423
rect 1460 1397 1486 1423
rect -123 1356 -97 1382
rect -33 1356 -7 1382
rect 143 1355 169 1381
rect 233 1355 259 1381
rect 773 1370 799 1396
rect -189 1325 -163 1351
rect 399 1335 425 1361
rect 859 1340 885 1366
rect 1045 1349 1071 1375
rect 1311 1348 1337 1374
rect -119 1278 -93 1304
rect -29 1278 -3 1304
rect 147 1277 173 1303
rect 237 1277 263 1303
rect 354 1274 380 1300
rect 390 1266 416 1292
rect 799 1268 825 1294
rect 859 1288 885 1314
rect 945 1295 971 1321
rect 1100 1308 1126 1334
rect 1190 1308 1216 1334
rect 1366 1307 1392 1333
rect 1456 1307 1482 1333
rect -178 1229 -152 1255
rect -119 1226 -93 1252
rect -29 1226 -3 1252
rect 88 1228 114 1254
rect 147 1225 173 1251
rect 237 1225 263 1251
rect 354 1222 380 1248
rect 859 1245 885 1271
rect 945 1243 971 1269
rect 1100 1256 1126 1282
rect 1190 1256 1216 1282
rect 1366 1255 1392 1281
rect 1456 1255 1482 1281
rect 1034 1225 1060 1251
rect -178 1177 -152 1203
rect 88 1176 114 1202
rect 313 1177 339 1203
rect 859 1193 885 1219
rect 1104 1178 1130 1204
rect 1194 1178 1220 1204
rect 1370 1177 1396 1203
rect 1460 1177 1486 1203
rect -123 1136 -97 1162
rect -33 1136 -7 1162
rect 143 1135 169 1161
rect 233 1135 259 1161
rect 399 1147 425 1173
rect 773 1137 799 1163
rect -123 1084 -97 1110
rect -33 1084 -7 1110
rect 143 1083 169 1109
rect 233 1083 259 1109
rect -189 1053 -163 1079
rect 339 1075 365 1101
rect 399 1095 425 1121
rect 485 1102 511 1128
rect 859 1107 885 1133
rect 1045 1129 1071 1155
rect 1104 1126 1130 1152
rect 1194 1126 1220 1152
rect 1311 1128 1337 1154
rect 1370 1125 1396 1151
rect 1460 1125 1486 1151
rect 399 1052 425 1078
rect 485 1050 511 1076
rect -119 1006 -93 1032
rect -29 1006 -3 1032
rect 147 1005 173 1031
rect 237 1005 263 1031
rect 399 1000 425 1026
rect 535 1017 561 1043
rect 573 1017 599 1043
rect 611 1017 637 1043
rect 649 1017 675 1043
rect 718 1018 744 1044
rect 799 1035 825 1061
rect 859 1055 885 1081
rect 945 1062 971 1088
rect 1045 1077 1071 1103
rect 1311 1076 1337 1102
rect 859 1012 885 1038
rect 1100 1036 1126 1062
rect 1190 1036 1216 1062
rect 945 1010 971 1036
rect 1366 1035 1392 1061
rect 1456 1035 1482 1061
rect -178 957 -152 983
rect -119 954 -93 980
rect -29 954 -3 980
rect 88 956 114 982
rect 147 953 173 979
rect 237 953 263 979
rect 354 939 380 965
rect 718 961 744 987
rect 859 960 885 986
rect 1100 984 1126 1010
rect 1190 984 1216 1010
rect 1366 983 1392 1009
rect 1456 983 1482 1009
rect 390 931 416 957
rect 1034 953 1060 979
rect -178 905 -152 931
rect 88 904 114 930
rect -123 864 -97 890
rect -33 864 -7 890
rect 143 863 169 889
rect 233 863 259 889
rect 354 887 380 913
rect 718 904 744 930
rect 773 904 799 930
rect 1104 906 1130 932
rect 1194 906 1220 932
rect 1370 905 1396 931
rect 1460 905 1486 931
rect 859 874 885 900
rect 313 842 339 868
rect 718 847 744 873
rect 1045 857 1071 883
rect -123 812 -97 838
rect -33 812 -7 838
rect 143 811 169 837
rect 233 811 259 837
rect 399 812 425 838
rect -189 781 -163 807
rect 799 802 825 828
rect 859 822 885 848
rect 945 829 971 855
rect 1104 854 1130 880
rect 1194 854 1220 880
rect 1311 856 1337 882
rect 1370 853 1396 879
rect 1460 853 1486 879
rect 1045 805 1071 831
rect -119 734 -93 760
rect -29 734 -3 760
rect 147 733 173 759
rect 237 733 263 759
rect 339 740 365 766
rect 399 760 425 786
rect 485 767 511 793
rect 859 779 885 805
rect 1311 804 1337 830
rect 945 777 971 803
rect 1100 764 1126 790
rect 1190 764 1216 790
rect 1366 763 1392 789
rect 1456 763 1482 789
rect 399 717 425 743
rect 485 715 511 741
rect 859 727 885 753
rect 1100 712 1126 738
rect 1190 712 1216 738
rect 1366 711 1392 737
rect 1456 711 1482 737
rect -178 685 -152 711
rect -119 682 -93 708
rect -29 682 -3 708
rect 88 684 114 710
rect 147 681 173 707
rect 237 681 263 707
rect 399 665 425 691
rect 773 671 799 697
rect 1034 681 1060 707
rect -178 633 -152 659
rect 88 632 114 658
rect 859 641 885 667
rect 1104 634 1130 660
rect 1194 634 1220 660
rect 1370 633 1396 659
rect 1460 633 1486 659
rect -123 592 -97 618
rect -33 592 -7 618
rect 143 591 169 617
rect 233 591 259 617
rect 354 604 380 630
rect 390 596 416 622
rect -123 540 -97 566
rect -33 540 -7 566
rect 143 539 169 565
rect 233 539 259 565
rect 354 552 380 578
rect 799 569 825 595
rect 859 589 885 615
rect 945 596 971 622
rect 1045 585 1071 611
rect 1104 582 1130 608
rect 1194 582 1220 608
rect 1311 584 1337 610
rect 1370 581 1396 607
rect 1460 581 1486 607
rect 859 546 885 572
rect 945 544 971 570
rect -189 509 -163 535
rect 1045 533 1071 559
rect 313 507 339 533
rect 1311 532 1337 558
rect -119 462 -93 488
rect -29 462 -3 488
rect 147 461 173 487
rect 237 461 263 487
rect 399 477 425 503
rect 859 494 885 520
rect 1100 492 1126 518
rect 1190 492 1216 518
rect 1366 491 1392 517
rect 1456 491 1482 517
rect -178 413 -152 439
rect -119 410 -93 436
rect -29 410 -3 436
rect 88 412 114 438
rect 147 409 173 435
rect 237 409 263 435
rect 339 405 365 431
rect 399 425 425 451
rect 485 432 511 458
rect 1100 440 1126 466
rect 1190 440 1216 466
rect 1366 439 1392 465
rect 1456 439 1482 465
rect 1034 409 1060 435
rect -178 361 -152 387
rect 88 360 114 386
rect 399 382 425 408
rect 485 380 511 406
rect 1104 362 1130 388
rect 1194 362 1220 388
rect 1370 361 1396 387
rect 1460 361 1486 387
rect -123 320 -97 346
rect -33 320 -7 346
rect 143 319 169 345
rect 233 319 259 345
rect 399 330 425 356
rect 1045 313 1071 339
rect 1104 310 1130 336
rect 1194 310 1220 336
rect 1311 312 1337 338
rect 1370 309 1396 335
rect 1460 309 1486 335
rect -123 268 -97 294
rect -33 268 -7 294
rect 143 267 169 293
rect 233 267 259 293
rect 354 269 380 295
rect -189 237 -163 263
rect 390 261 416 287
rect 1045 261 1071 287
rect 1311 260 1337 286
rect 354 217 380 243
rect -119 190 -93 216
rect -29 190 -3 216
rect 147 189 173 215
rect 237 189 263 215
rect -178 141 -152 167
rect -119 138 -93 164
rect -29 138 -3 164
rect 88 140 114 166
rect 147 137 173 163
rect 237 137 263 163
rect -178 89 -152 115
rect 88 88 114 114
rect -123 48 -97 74
rect -33 48 -7 74
rect 143 47 169 73
rect 233 47 259 73
rect -123 -4 -97 22
rect -33 -4 -7 22
rect 143 -5 169 21
rect 233 -5 259 21
rect -189 -35 -163 -9
rect -119 -82 -93 -56
rect -29 -82 -3 -56
rect 147 -83 173 -57
rect 237 -83 263 -57
rect -178 -131 -152 -105
rect -119 -134 -93 -108
rect -29 -134 -3 -108
rect 88 -132 114 -106
rect 147 -135 173 -109
rect 237 -135 263 -109
rect -178 -183 -152 -157
rect 88 -184 114 -158
<< ntransistor >>
rect -163 1946 -155 1948
rect -73 1946 -65 1948
rect 103 1945 111 1947
rect 193 1945 201 1947
rect -141 1938 -133 1940
rect -51 1938 -43 1940
rect 125 1937 133 1939
rect 215 1937 223 1939
rect -177 1855 -175 1863
rect -159 1816 -151 1818
rect -69 1816 -61 1818
rect 107 1815 115 1817
rect 197 1815 205 1817
rect -137 1808 -129 1810
rect -47 1808 -39 1810
rect 129 1807 137 1809
rect 219 1807 227 1809
rect -218 1767 -210 1769
rect 48 1766 56 1768
rect -196 1759 -188 1761
rect 70 1758 78 1760
rect -163 1674 -155 1676
rect -73 1674 -65 1676
rect 103 1673 111 1675
rect 193 1673 201 1675
rect -141 1666 -133 1668
rect -51 1666 -43 1668
rect 125 1665 133 1667
rect 215 1665 223 1667
rect -177 1583 -175 1591
rect 1060 1574 1068 1576
rect 1150 1574 1158 1576
rect 1326 1573 1334 1575
rect 1416 1573 1424 1575
rect 1082 1566 1090 1568
rect 1172 1566 1180 1568
rect 1348 1565 1356 1567
rect 1438 1565 1446 1567
rect -159 1544 -151 1546
rect -69 1544 -61 1546
rect 107 1543 115 1545
rect 197 1543 205 1545
rect -137 1536 -129 1538
rect -47 1536 -39 1538
rect 129 1535 137 1537
rect 219 1535 227 1537
rect -218 1495 -210 1497
rect 325 1498 327 1506
rect 48 1494 56 1496
rect -196 1487 -188 1489
rect 70 1486 78 1488
rect 1046 1483 1048 1491
rect 359 1476 367 1478
rect 381 1468 389 1470
rect 1064 1444 1072 1446
rect 1154 1444 1162 1446
rect 1330 1443 1338 1445
rect 1420 1443 1428 1445
rect 1086 1436 1094 1438
rect 1176 1436 1184 1438
rect 445 1431 453 1433
rect 1352 1435 1360 1437
rect 1442 1435 1450 1437
rect 325 1422 333 1424
rect 467 1423 475 1425
rect -163 1402 -155 1404
rect -73 1402 -65 1404
rect 103 1401 111 1403
rect 193 1401 201 1403
rect -141 1394 -133 1396
rect -51 1394 -43 1396
rect 125 1393 133 1395
rect 215 1393 223 1395
rect 1005 1395 1013 1397
rect 1271 1394 1279 1396
rect 1027 1387 1035 1389
rect 359 1381 367 1383
rect 1293 1386 1301 1388
rect 381 1373 389 1375
rect 785 1356 787 1364
rect 819 1334 827 1336
rect 841 1326 849 1328
rect -177 1311 -175 1319
rect 1060 1302 1068 1304
rect 1150 1302 1158 1304
rect 1326 1301 1334 1303
rect 1416 1301 1424 1303
rect 1082 1294 1090 1296
rect 1172 1294 1180 1296
rect 905 1289 913 1291
rect 1348 1293 1356 1295
rect 1438 1293 1446 1295
rect 785 1280 793 1282
rect 927 1281 935 1283
rect -159 1272 -151 1274
rect -69 1272 -61 1274
rect 107 1271 115 1273
rect 197 1271 205 1273
rect 314 1268 322 1270
rect -137 1264 -129 1266
rect -47 1264 -39 1266
rect 129 1263 137 1265
rect 219 1263 227 1265
rect 336 1260 344 1262
rect 402 1252 404 1260
rect 819 1239 827 1241
rect -218 1223 -210 1225
rect 841 1231 849 1233
rect 48 1222 56 1224
rect -196 1215 -188 1217
rect 70 1214 78 1216
rect 1046 1211 1048 1219
rect 1064 1172 1072 1174
rect 1154 1172 1162 1174
rect 1330 1171 1338 1173
rect 1420 1171 1428 1173
rect 325 1163 327 1171
rect 1086 1164 1094 1166
rect 1176 1164 1184 1166
rect 1352 1163 1360 1165
rect 1442 1163 1450 1165
rect 359 1141 367 1143
rect -163 1130 -155 1132
rect -73 1130 -65 1132
rect 381 1133 389 1135
rect 103 1129 111 1131
rect 193 1129 201 1131
rect -141 1122 -133 1124
rect -51 1122 -43 1124
rect 125 1121 133 1123
rect 215 1121 223 1123
rect 785 1123 787 1131
rect 1005 1123 1013 1125
rect 1271 1122 1279 1124
rect 1027 1115 1035 1117
rect 1293 1114 1301 1116
rect 819 1101 827 1103
rect 445 1096 453 1098
rect 841 1093 849 1095
rect 325 1087 333 1089
rect 467 1088 475 1090
rect 905 1056 913 1058
rect -177 1039 -175 1047
rect 359 1046 367 1048
rect 785 1047 793 1049
rect 927 1048 935 1050
rect 381 1038 389 1040
rect 1060 1030 1068 1032
rect 1150 1030 1158 1032
rect 1326 1029 1334 1031
rect 1416 1029 1424 1031
rect -159 1000 -151 1002
rect -69 1000 -61 1002
rect 1082 1022 1090 1024
rect 1172 1022 1180 1024
rect 730 1004 732 1012
rect 1348 1021 1356 1023
rect 1438 1021 1446 1023
rect 819 1006 827 1008
rect 107 999 115 1001
rect 197 999 205 1001
rect 841 998 849 1000
rect -137 992 -129 994
rect -47 992 -39 994
rect 129 991 137 993
rect 219 991 227 993
rect 661 983 663 991
rect 691 984 693 992
rect -218 951 -210 953
rect 653 953 655 961
rect 48 950 56 952
rect -196 943 -188 945
rect 70 942 78 944
rect 623 942 625 950
rect 730 947 732 955
rect 1046 939 1048 947
rect 314 933 322 935
rect 336 925 344 927
rect 402 917 404 925
rect 615 912 617 920
rect 585 901 587 909
rect 1064 900 1072 902
rect 1154 900 1162 902
rect 1330 899 1338 901
rect 1420 899 1428 901
rect 730 890 732 898
rect 785 890 787 898
rect 1086 892 1094 894
rect 1176 892 1184 894
rect 1352 891 1360 893
rect 1442 891 1450 893
rect 577 871 579 879
rect 819 868 827 870
rect -163 858 -155 860
rect -73 858 -65 860
rect 547 860 549 868
rect 103 857 111 859
rect 193 857 201 859
rect -141 850 -133 852
rect -51 850 -43 852
rect 125 849 133 851
rect 215 849 223 851
rect 841 860 849 862
rect 1005 851 1013 853
rect 1271 850 1279 852
rect 1027 843 1035 845
rect 325 828 327 836
rect 539 831 541 839
rect 730 833 732 841
rect 1293 842 1301 844
rect 905 823 913 825
rect 785 814 793 816
rect 927 815 935 817
rect 359 806 367 808
rect 531 802 533 810
rect 381 798 389 800
rect -177 767 -175 775
rect 819 773 827 775
rect 841 765 849 767
rect 445 761 453 763
rect 1060 758 1068 760
rect 1150 758 1158 760
rect 1326 757 1334 759
rect 1416 757 1424 759
rect 325 752 333 754
rect 467 753 475 755
rect 1082 750 1090 752
rect 1172 750 1180 752
rect 1348 749 1356 751
rect 1438 749 1446 751
rect -159 728 -151 730
rect -69 728 -61 730
rect 107 727 115 729
rect 197 727 205 729
rect -137 720 -129 722
rect -47 720 -39 722
rect 129 719 137 721
rect 219 719 227 721
rect 359 711 367 713
rect 381 703 389 705
rect -218 679 -210 681
rect 48 678 56 680
rect -196 671 -188 673
rect 70 670 78 672
rect 1046 667 1048 675
rect 785 657 787 665
rect 819 635 827 637
rect 841 627 849 629
rect 1064 628 1072 630
rect 1154 628 1162 630
rect 1330 627 1338 629
rect 1420 627 1428 629
rect 1086 620 1094 622
rect 1176 620 1184 622
rect 1352 619 1360 621
rect 1442 619 1450 621
rect 314 598 322 600
rect -163 586 -155 588
rect -73 586 -65 588
rect 336 590 344 592
rect 103 585 111 587
rect 193 585 201 587
rect 402 582 404 590
rect 905 590 913 592
rect -141 578 -133 580
rect -51 578 -43 580
rect 125 577 133 579
rect 215 577 223 579
rect 785 581 793 583
rect 927 582 935 584
rect 1005 579 1013 581
rect 1271 578 1279 580
rect 1027 571 1035 573
rect 1293 570 1301 572
rect 819 540 827 542
rect 841 532 849 534
rect -177 495 -175 503
rect 325 493 327 501
rect 1060 486 1068 488
rect 1150 486 1158 488
rect 1326 485 1334 487
rect 1416 485 1424 487
rect 1082 478 1090 480
rect 1172 478 1180 480
rect 359 471 367 473
rect 1348 477 1356 479
rect 1438 477 1446 479
rect 381 463 389 465
rect -159 456 -151 458
rect -69 456 -61 458
rect 107 455 115 457
rect 197 455 205 457
rect -137 448 -129 450
rect -47 448 -39 450
rect 129 447 137 449
rect 219 447 227 449
rect -218 407 -210 409
rect 445 426 453 428
rect 325 417 333 419
rect 467 418 475 420
rect 48 406 56 408
rect -196 399 -188 401
rect 70 398 78 400
rect 1046 395 1048 403
rect 359 376 367 378
rect 381 368 389 370
rect 1064 356 1072 358
rect 1154 356 1162 358
rect 1330 355 1338 357
rect 1420 355 1428 357
rect 1086 348 1094 350
rect 1176 348 1184 350
rect 1352 347 1360 349
rect 1442 347 1450 349
rect -163 314 -155 316
rect -73 314 -65 316
rect 103 313 111 315
rect 193 313 201 315
rect -141 306 -133 308
rect -51 306 -43 308
rect 1005 307 1013 309
rect 125 305 133 307
rect 215 305 223 307
rect 1271 306 1279 308
rect 1027 299 1035 301
rect 1293 298 1301 300
rect 314 263 322 265
rect 336 255 344 257
rect 402 247 404 255
rect -177 223 -175 231
rect -159 184 -151 186
rect -69 184 -61 186
rect 107 183 115 185
rect 197 183 205 185
rect -137 176 -129 178
rect -47 176 -39 178
rect 129 175 137 177
rect 219 175 227 177
rect -218 135 -210 137
rect 48 134 56 136
rect -196 127 -188 129
rect 70 126 78 128
rect -163 42 -155 44
rect -73 42 -65 44
rect 103 41 111 43
rect 193 41 201 43
rect -141 34 -133 36
rect -51 34 -43 36
rect 125 33 133 35
rect 215 33 223 35
rect -177 -49 -175 -41
rect -159 -88 -151 -86
rect -69 -88 -61 -86
rect 107 -89 115 -87
rect 197 -89 205 -87
rect -137 -96 -129 -94
rect -47 -96 -39 -94
rect 129 -97 137 -95
rect 219 -97 227 -95
rect -218 -137 -210 -135
rect 48 -138 56 -136
rect -196 -145 -188 -143
rect 70 -146 78 -144
<< ptransistor >>
rect -117 1964 -109 1966
rect -27 1964 -19 1966
rect 149 1963 157 1965
rect 239 1963 247 1965
rect -117 1912 -109 1914
rect -27 1912 -19 1914
rect 149 1911 157 1913
rect 239 1911 247 1913
rect -177 1875 -175 1883
rect -113 1834 -105 1836
rect -23 1834 -15 1836
rect 153 1833 161 1835
rect 243 1833 251 1835
rect -172 1785 -164 1787
rect 94 1784 102 1786
rect -113 1782 -105 1784
rect -23 1782 -15 1784
rect 153 1781 161 1783
rect 243 1781 251 1783
rect -172 1733 -164 1735
rect 94 1732 102 1734
rect -117 1692 -109 1694
rect -27 1692 -19 1694
rect 149 1691 157 1693
rect 239 1691 247 1693
rect -117 1640 -109 1642
rect -27 1640 -19 1642
rect 149 1639 157 1641
rect 239 1639 247 1641
rect -177 1603 -175 1611
rect 1106 1592 1114 1594
rect 1196 1592 1204 1594
rect 1372 1591 1380 1593
rect 1462 1591 1470 1593
rect -113 1562 -105 1564
rect -23 1562 -15 1564
rect 153 1561 161 1563
rect 243 1561 251 1563
rect 1106 1540 1114 1542
rect 1196 1540 1204 1542
rect 1372 1539 1380 1541
rect 1462 1539 1470 1541
rect -172 1513 -164 1515
rect 325 1518 327 1526
rect 94 1512 102 1514
rect -113 1510 -105 1512
rect -23 1510 -15 1512
rect 153 1509 161 1511
rect 243 1509 251 1511
rect 1046 1503 1048 1511
rect 405 1494 413 1496
rect -172 1461 -164 1463
rect 94 1460 102 1462
rect 1110 1462 1118 1464
rect 1200 1462 1208 1464
rect 1376 1461 1384 1463
rect 1466 1461 1474 1463
rect 491 1449 499 1451
rect 405 1442 413 1444
rect -117 1420 -109 1422
rect -27 1420 -19 1422
rect 345 1422 353 1424
rect 149 1419 157 1421
rect 239 1419 247 1421
rect 1051 1413 1059 1415
rect 1317 1412 1325 1414
rect 1110 1410 1118 1412
rect 1200 1410 1208 1412
rect 405 1399 413 1401
rect 491 1397 499 1399
rect 1376 1409 1384 1411
rect 1466 1409 1474 1411
rect 785 1376 787 1384
rect -117 1368 -109 1370
rect -27 1368 -19 1370
rect 149 1367 157 1369
rect 239 1367 247 1369
rect 1051 1361 1059 1363
rect 1317 1360 1325 1362
rect 865 1352 873 1354
rect 405 1347 413 1349
rect -177 1331 -175 1339
rect 1106 1320 1114 1322
rect 1196 1320 1204 1322
rect 1372 1319 1380 1321
rect 1462 1319 1470 1321
rect 951 1307 959 1309
rect 865 1300 873 1302
rect -113 1290 -105 1292
rect -23 1290 -15 1292
rect 153 1289 161 1291
rect 243 1289 251 1291
rect 360 1286 368 1288
rect 805 1280 813 1282
rect 402 1272 404 1280
rect 1106 1268 1114 1270
rect 1196 1268 1204 1270
rect 865 1257 873 1259
rect 1372 1267 1380 1269
rect 1462 1267 1470 1269
rect 951 1255 959 1257
rect -172 1241 -164 1243
rect 94 1240 102 1242
rect -113 1238 -105 1240
rect -23 1238 -15 1240
rect 153 1237 161 1239
rect 243 1237 251 1239
rect 360 1234 368 1236
rect 1046 1231 1048 1239
rect 865 1205 873 1207
rect -172 1189 -164 1191
rect 94 1188 102 1190
rect 325 1183 327 1191
rect 1110 1190 1118 1192
rect 1200 1190 1208 1192
rect 1376 1189 1384 1191
rect 1466 1189 1474 1191
rect 405 1159 413 1161
rect -117 1148 -109 1150
rect -27 1148 -19 1150
rect 149 1147 157 1149
rect 239 1147 247 1149
rect 785 1143 787 1151
rect 1051 1141 1059 1143
rect 1317 1140 1325 1142
rect 1110 1138 1118 1140
rect 1200 1138 1208 1140
rect 1376 1137 1384 1139
rect 1466 1137 1474 1139
rect 865 1119 873 1121
rect 491 1114 499 1116
rect 405 1107 413 1109
rect -117 1096 -109 1098
rect -27 1096 -19 1098
rect 149 1095 157 1097
rect 239 1095 247 1097
rect 345 1087 353 1089
rect 1051 1089 1059 1091
rect 1317 1088 1325 1090
rect 951 1074 959 1076
rect -177 1059 -175 1067
rect 405 1064 413 1066
rect 865 1067 873 1069
rect 491 1062 499 1064
rect 805 1047 813 1049
rect 1106 1048 1114 1050
rect 1196 1048 1204 1050
rect 1372 1047 1380 1049
rect 1462 1047 1470 1049
rect -113 1018 -105 1020
rect -23 1018 -15 1020
rect 547 1023 549 1031
rect 585 1023 587 1031
rect 623 1023 625 1031
rect 661 1023 663 1031
rect 730 1024 732 1032
rect 865 1024 873 1026
rect 153 1017 161 1019
rect 243 1017 251 1019
rect 405 1012 413 1014
rect 951 1022 959 1024
rect 1106 996 1114 998
rect 1196 996 1204 998
rect 1372 995 1380 997
rect 1462 995 1470 997
rect -172 969 -164 971
rect 94 968 102 970
rect -113 966 -105 968
rect -23 966 -15 968
rect 153 965 161 967
rect 243 965 251 967
rect 730 967 732 975
rect 865 972 873 974
rect 1046 959 1048 967
rect 360 951 368 953
rect 402 937 404 945
rect -172 917 -164 919
rect 94 916 102 918
rect 1110 918 1118 920
rect 1200 918 1208 920
rect 730 910 732 918
rect 785 910 787 918
rect 1376 917 1384 919
rect 1466 917 1474 919
rect 360 899 368 901
rect -117 876 -109 878
rect -27 876 -19 878
rect 865 886 873 888
rect 149 875 157 877
rect 239 875 247 877
rect 1051 869 1059 871
rect 1317 868 1325 870
rect 1110 866 1118 868
rect 1200 866 1208 868
rect 325 848 327 856
rect 730 853 732 861
rect 1376 865 1384 867
rect 1466 865 1474 867
rect 951 841 959 843
rect -117 824 -109 826
rect -27 824 -19 826
rect 865 834 873 836
rect 149 823 157 825
rect 239 823 247 825
rect 405 824 413 826
rect 1051 817 1059 819
rect 805 814 813 816
rect 1317 816 1325 818
rect -177 787 -175 795
rect 865 791 873 793
rect 951 789 959 791
rect 491 779 499 781
rect 1106 776 1114 778
rect 1196 776 1204 778
rect 405 772 413 774
rect 1372 775 1380 777
rect 1462 775 1470 777
rect -113 746 -105 748
rect -23 746 -15 748
rect 345 752 353 754
rect 153 745 161 747
rect 243 745 251 747
rect 865 739 873 741
rect 405 729 413 731
rect 491 727 499 729
rect 1106 724 1114 726
rect 1196 724 1204 726
rect 1372 723 1380 725
rect 1462 723 1470 725
rect -172 697 -164 699
rect 94 696 102 698
rect -113 694 -105 696
rect -23 694 -15 696
rect 153 693 161 695
rect 243 693 251 695
rect 1046 687 1048 695
rect 405 677 413 679
rect 785 677 787 685
rect 865 653 873 655
rect -172 645 -164 647
rect 94 644 102 646
rect 1110 646 1118 648
rect 1200 646 1208 648
rect 1376 645 1384 647
rect 1466 645 1474 647
rect 360 616 368 618
rect -117 604 -109 606
rect -27 604 -19 606
rect 149 603 157 605
rect 239 603 247 605
rect 402 602 404 610
rect 951 608 959 610
rect 865 601 873 603
rect 1051 597 1059 599
rect 1317 596 1325 598
rect 1110 594 1118 596
rect 1200 594 1208 596
rect 805 581 813 583
rect 1376 593 1384 595
rect 1466 593 1474 595
rect 360 564 368 566
rect -117 552 -109 554
rect -27 552 -19 554
rect 865 558 873 560
rect 951 556 959 558
rect 149 551 157 553
rect 239 551 247 553
rect 1051 545 1059 547
rect 1317 544 1325 546
rect -177 515 -175 523
rect 325 513 327 521
rect 865 506 873 508
rect 1106 504 1114 506
rect 1196 504 1204 506
rect 1372 503 1380 505
rect 1462 503 1470 505
rect 405 489 413 491
rect -113 474 -105 476
rect -23 474 -15 476
rect 153 473 161 475
rect 243 473 251 475
rect 1106 452 1114 454
rect 1196 452 1204 454
rect 491 444 499 446
rect 1372 451 1380 453
rect 1462 451 1470 453
rect 405 437 413 439
rect -172 425 -164 427
rect 94 424 102 426
rect -113 422 -105 424
rect -23 422 -15 424
rect 153 421 161 423
rect 243 421 251 423
rect 345 417 353 419
rect 1046 415 1048 423
rect 405 394 413 396
rect 491 392 499 394
rect -172 373 -164 375
rect 94 372 102 374
rect 1110 374 1118 376
rect 1200 374 1208 376
rect 1376 373 1384 375
rect 1466 373 1474 375
rect 405 342 413 344
rect -117 332 -109 334
rect -27 332 -19 334
rect 149 331 157 333
rect 239 331 247 333
rect 1051 325 1059 327
rect 1317 324 1325 326
rect 1110 322 1118 324
rect 1200 322 1208 324
rect 1376 321 1384 323
rect 1466 321 1474 323
rect -117 280 -109 282
rect -27 280 -19 282
rect 360 281 368 283
rect 149 279 157 281
rect 239 279 247 281
rect 402 267 404 275
rect 1051 273 1059 275
rect 1317 272 1325 274
rect -177 243 -175 251
rect 360 229 368 231
rect -113 202 -105 204
rect -23 202 -15 204
rect 153 201 161 203
rect 243 201 251 203
rect -172 153 -164 155
rect 94 152 102 154
rect -113 150 -105 152
rect -23 150 -15 152
rect 153 149 161 151
rect 243 149 251 151
rect -172 101 -164 103
rect 94 100 102 102
rect -117 60 -109 62
rect -27 60 -19 62
rect 149 59 157 61
rect 239 59 247 61
rect -117 8 -109 10
rect -27 8 -19 10
rect 149 7 157 9
rect 239 7 247 9
rect -177 -29 -175 -21
rect -113 -70 -105 -68
rect -23 -70 -15 -68
rect 153 -71 161 -69
rect 243 -71 251 -69
rect -172 -119 -164 -117
rect 94 -120 102 -118
rect -113 -122 -105 -120
rect -23 -122 -15 -120
rect 153 -123 161 -121
rect 243 -123 251 -121
rect -172 -171 -164 -169
rect 94 -172 102 -170
<< ndiffusion >>
rect -163 1948 -155 1949
rect -73 1948 -65 1949
rect 103 1947 111 1948
rect 193 1947 201 1948
rect -163 1945 -155 1946
rect -73 1945 -65 1946
rect -141 1940 -133 1941
rect -51 1940 -43 1941
rect 103 1944 111 1945
rect 193 1944 201 1945
rect 125 1939 133 1940
rect 215 1939 223 1940
rect -141 1937 -133 1938
rect -51 1937 -43 1938
rect 125 1936 133 1937
rect 215 1936 223 1937
rect -178 1855 -177 1863
rect -175 1855 -174 1863
rect -159 1818 -151 1819
rect -69 1818 -61 1819
rect 107 1817 115 1818
rect 197 1817 205 1818
rect -159 1815 -151 1816
rect -69 1815 -61 1816
rect -137 1810 -129 1811
rect -47 1810 -39 1811
rect 107 1814 115 1815
rect 197 1814 205 1815
rect 129 1809 137 1810
rect 219 1809 227 1810
rect -137 1807 -129 1808
rect -47 1807 -39 1808
rect 129 1806 137 1807
rect 219 1806 227 1807
rect -218 1769 -210 1770
rect 48 1768 56 1769
rect -218 1766 -210 1767
rect -196 1761 -188 1762
rect 48 1765 56 1766
rect 70 1760 78 1761
rect -196 1758 -188 1759
rect 70 1757 78 1758
rect -163 1676 -155 1677
rect -73 1676 -65 1677
rect 103 1675 111 1676
rect 193 1675 201 1676
rect -163 1673 -155 1674
rect -73 1673 -65 1674
rect -141 1668 -133 1669
rect -51 1668 -43 1669
rect 103 1672 111 1673
rect 193 1672 201 1673
rect 125 1667 133 1668
rect 215 1667 223 1668
rect -141 1665 -133 1666
rect -51 1665 -43 1666
rect 125 1664 133 1665
rect 215 1664 223 1665
rect -178 1583 -177 1591
rect -175 1583 -174 1591
rect 1060 1576 1068 1577
rect 1150 1576 1158 1577
rect 1326 1575 1334 1576
rect 1416 1575 1424 1576
rect 1060 1573 1068 1574
rect 1150 1573 1158 1574
rect 1082 1568 1090 1569
rect 1172 1568 1180 1569
rect 1326 1572 1334 1573
rect 1416 1572 1424 1573
rect 1348 1567 1356 1568
rect 1438 1567 1446 1568
rect 1082 1565 1090 1566
rect 1172 1565 1180 1566
rect -159 1546 -151 1547
rect -69 1546 -61 1547
rect 1348 1564 1356 1565
rect 1438 1564 1446 1565
rect 107 1545 115 1546
rect 197 1545 205 1546
rect -159 1543 -151 1544
rect -69 1543 -61 1544
rect -137 1538 -129 1539
rect -47 1538 -39 1539
rect 107 1542 115 1543
rect 197 1542 205 1543
rect 129 1537 137 1538
rect 219 1537 227 1538
rect -137 1535 -129 1536
rect -47 1535 -39 1536
rect 129 1534 137 1535
rect 219 1534 227 1535
rect -218 1497 -210 1498
rect 48 1496 56 1497
rect 324 1498 325 1506
rect 327 1498 328 1506
rect -218 1494 -210 1495
rect -196 1489 -188 1490
rect 48 1493 56 1494
rect 70 1488 78 1489
rect -196 1486 -188 1487
rect 70 1485 78 1486
rect 359 1478 367 1479
rect 1045 1483 1046 1491
rect 1048 1483 1049 1491
rect 359 1475 367 1476
rect 381 1470 389 1471
rect 381 1467 389 1468
rect 1064 1446 1072 1447
rect 1154 1446 1162 1447
rect 1330 1445 1338 1446
rect 1420 1445 1428 1446
rect 1064 1443 1072 1444
rect 1154 1443 1162 1444
rect 445 1433 453 1434
rect 1086 1438 1094 1439
rect 1176 1438 1184 1439
rect 1330 1442 1338 1443
rect 1420 1442 1428 1443
rect 1352 1437 1360 1438
rect 1442 1437 1450 1438
rect 325 1424 333 1425
rect 445 1430 453 1431
rect 1086 1435 1094 1436
rect 1176 1435 1184 1436
rect 467 1425 475 1426
rect 1352 1434 1360 1435
rect 1442 1434 1450 1435
rect 325 1421 333 1422
rect 467 1422 475 1423
rect -163 1404 -155 1405
rect -73 1404 -65 1405
rect 103 1403 111 1404
rect 193 1403 201 1404
rect -163 1401 -155 1402
rect -73 1401 -65 1402
rect -141 1396 -133 1397
rect -51 1396 -43 1397
rect 103 1400 111 1401
rect 193 1400 201 1401
rect 125 1395 133 1396
rect 215 1395 223 1396
rect -141 1393 -133 1394
rect -51 1393 -43 1394
rect 1005 1397 1013 1398
rect 125 1392 133 1393
rect 215 1392 223 1393
rect 1271 1396 1279 1397
rect 1005 1394 1013 1395
rect 1027 1389 1035 1390
rect 1271 1393 1279 1394
rect 359 1383 367 1384
rect 1293 1388 1301 1389
rect 359 1380 367 1381
rect 1027 1386 1035 1387
rect 381 1375 389 1376
rect 381 1372 389 1373
rect 1293 1385 1301 1386
rect 784 1356 785 1364
rect 787 1356 788 1364
rect 819 1336 827 1337
rect 819 1333 827 1334
rect 841 1328 849 1329
rect -178 1311 -177 1319
rect -175 1311 -174 1319
rect 841 1325 849 1326
rect 1060 1304 1068 1305
rect 1150 1304 1158 1305
rect 1326 1303 1334 1304
rect 1416 1303 1424 1304
rect 1060 1301 1068 1302
rect 1150 1301 1158 1302
rect 905 1291 913 1292
rect 1082 1296 1090 1297
rect 1172 1296 1180 1297
rect 1326 1300 1334 1301
rect 1416 1300 1424 1301
rect 1348 1295 1356 1296
rect 1438 1295 1446 1296
rect -159 1274 -151 1275
rect -69 1274 -61 1275
rect 785 1282 793 1283
rect 905 1288 913 1289
rect 1082 1293 1090 1294
rect 1172 1293 1180 1294
rect 927 1283 935 1284
rect 1348 1292 1356 1293
rect 1438 1292 1446 1293
rect 107 1273 115 1274
rect 197 1273 205 1274
rect -159 1271 -151 1272
rect -69 1271 -61 1272
rect -137 1266 -129 1267
rect -47 1266 -39 1267
rect 107 1270 115 1271
rect 197 1270 205 1271
rect 314 1270 322 1271
rect 785 1279 793 1280
rect 927 1280 935 1281
rect 129 1265 137 1266
rect 219 1265 227 1266
rect 314 1267 322 1268
rect -137 1263 -129 1264
rect -47 1263 -39 1264
rect 129 1262 137 1263
rect 219 1262 227 1263
rect 336 1262 344 1263
rect 336 1259 344 1260
rect 401 1252 402 1260
rect 404 1252 405 1260
rect 819 1241 827 1242
rect -218 1225 -210 1226
rect 48 1224 56 1225
rect 819 1238 827 1239
rect 841 1233 849 1234
rect -218 1222 -210 1223
rect 841 1230 849 1231
rect -196 1217 -188 1218
rect 48 1221 56 1222
rect 70 1216 78 1217
rect -196 1214 -188 1215
rect 70 1213 78 1214
rect 1045 1211 1046 1219
rect 1048 1211 1049 1219
rect 1064 1174 1072 1175
rect 1154 1174 1162 1175
rect 1330 1173 1338 1174
rect 1420 1173 1428 1174
rect 1064 1171 1072 1172
rect 1154 1171 1162 1172
rect 324 1163 325 1171
rect 327 1163 328 1171
rect 1086 1166 1094 1167
rect 1176 1166 1184 1167
rect 1330 1170 1338 1171
rect 1420 1170 1428 1171
rect 1352 1165 1360 1166
rect 1442 1165 1450 1166
rect 1086 1163 1094 1164
rect 1176 1163 1184 1164
rect 1352 1162 1360 1163
rect 1442 1162 1450 1163
rect 359 1143 367 1144
rect -163 1132 -155 1133
rect -73 1132 -65 1133
rect 359 1140 367 1141
rect 103 1131 111 1132
rect 193 1131 201 1132
rect 381 1135 389 1136
rect -163 1129 -155 1130
rect -73 1129 -65 1130
rect -141 1124 -133 1125
rect -51 1124 -43 1125
rect 103 1128 111 1129
rect 193 1128 201 1129
rect 381 1132 389 1133
rect 125 1123 133 1124
rect 215 1123 223 1124
rect -141 1121 -133 1122
rect -51 1121 -43 1122
rect 125 1120 133 1121
rect 215 1120 223 1121
rect 784 1123 785 1131
rect 787 1123 788 1131
rect 1005 1125 1013 1126
rect 1271 1124 1279 1125
rect 1005 1122 1013 1123
rect 1027 1117 1035 1118
rect 1271 1121 1279 1122
rect 1293 1116 1301 1117
rect 445 1098 453 1099
rect 819 1103 827 1104
rect 1027 1114 1035 1115
rect 1293 1113 1301 1114
rect 819 1100 827 1101
rect 325 1089 333 1090
rect 445 1095 453 1096
rect 841 1095 849 1096
rect 467 1090 475 1091
rect 325 1086 333 1087
rect 467 1087 475 1088
rect 841 1092 849 1093
rect 905 1058 913 1059
rect 359 1048 367 1049
rect 785 1049 793 1050
rect 905 1055 913 1056
rect 927 1050 935 1051
rect -178 1039 -177 1047
rect -175 1039 -174 1047
rect 785 1046 793 1047
rect 359 1045 367 1046
rect 381 1040 389 1041
rect 927 1047 935 1048
rect 381 1037 389 1038
rect 1060 1032 1068 1033
rect 1150 1032 1158 1033
rect 1326 1031 1334 1032
rect 1416 1031 1424 1032
rect 1060 1029 1068 1030
rect 1150 1029 1158 1030
rect 1082 1024 1090 1025
rect 1172 1024 1180 1025
rect 1326 1028 1334 1029
rect 1416 1028 1424 1029
rect -159 1002 -151 1003
rect -69 1002 -61 1003
rect 107 1001 115 1002
rect 197 1001 205 1002
rect 1348 1023 1356 1024
rect 1438 1023 1446 1024
rect 729 1004 730 1012
rect 732 1004 733 1012
rect 819 1008 827 1009
rect 1082 1021 1090 1022
rect 1172 1021 1180 1022
rect 1348 1020 1356 1021
rect 1438 1020 1446 1021
rect 819 1005 827 1006
rect -159 999 -151 1000
rect -69 999 -61 1000
rect 841 1000 849 1001
rect -137 994 -129 995
rect -47 994 -39 995
rect 107 998 115 999
rect 197 998 205 999
rect 129 993 137 994
rect 219 993 227 994
rect -137 991 -129 992
rect -47 991 -39 992
rect 129 990 137 991
rect 219 990 227 991
rect 660 983 661 991
rect 663 983 664 991
rect 690 984 691 992
rect 693 984 694 992
rect 841 997 849 998
rect -218 953 -210 954
rect 48 952 56 953
rect 652 953 653 961
rect 655 953 656 961
rect -218 950 -210 951
rect -196 945 -188 946
rect 48 949 56 950
rect 70 944 78 945
rect -196 942 -188 943
rect 70 941 78 942
rect 314 935 322 936
rect 622 942 623 950
rect 625 942 626 950
rect 729 947 730 955
rect 732 947 733 955
rect 1045 939 1046 947
rect 1048 939 1049 947
rect 314 932 322 933
rect 336 927 344 928
rect 336 924 344 925
rect 401 917 402 925
rect 404 917 405 925
rect 614 912 615 920
rect 617 912 618 920
rect 584 901 585 909
rect 587 901 588 909
rect 1064 902 1072 903
rect 1154 902 1162 903
rect 1330 901 1338 902
rect 1420 901 1428 902
rect 1064 899 1072 900
rect 1154 899 1162 900
rect 729 890 730 898
rect 732 890 733 898
rect 784 890 785 898
rect 787 890 788 898
rect 1086 894 1094 895
rect 1176 894 1184 895
rect 1330 898 1338 899
rect 1420 898 1428 899
rect 1352 893 1360 894
rect 1442 893 1450 894
rect 1086 891 1094 892
rect 1176 891 1184 892
rect -163 860 -155 861
rect -73 860 -65 861
rect 576 871 577 879
rect 579 871 580 879
rect 1352 890 1360 891
rect 1442 890 1450 891
rect 819 870 827 871
rect 103 859 111 860
rect 193 859 201 860
rect 546 860 547 868
rect 549 860 550 868
rect 819 867 827 868
rect 841 862 849 863
rect -163 857 -155 858
rect -73 857 -65 858
rect -141 852 -133 853
rect -51 852 -43 853
rect 103 856 111 857
rect 193 856 201 857
rect 125 851 133 852
rect 215 851 223 852
rect -141 849 -133 850
rect -51 849 -43 850
rect 125 848 133 849
rect 215 848 223 849
rect 841 859 849 860
rect 1005 853 1013 854
rect 1271 852 1279 853
rect 1005 850 1013 851
rect 1027 845 1035 846
rect 1271 849 1279 850
rect 1293 844 1301 845
rect 324 828 325 836
rect 327 828 328 836
rect 538 831 539 839
rect 541 831 542 839
rect 729 833 730 841
rect 732 833 733 841
rect 1027 842 1035 843
rect 905 825 913 826
rect 1293 841 1301 842
rect 785 816 793 817
rect 905 822 913 823
rect 927 817 935 818
rect 359 808 367 809
rect 785 813 793 814
rect 359 805 367 806
rect 530 802 531 810
rect 533 802 534 810
rect 927 814 935 815
rect 381 800 389 801
rect 381 797 389 798
rect -178 767 -177 775
rect -175 767 -174 775
rect 819 775 827 776
rect 819 772 827 773
rect 445 763 453 764
rect 841 767 849 768
rect 325 754 333 755
rect 445 760 453 761
rect 841 764 849 765
rect 1060 760 1068 761
rect 1150 760 1158 761
rect 1326 759 1334 760
rect 1416 759 1424 760
rect 1060 757 1068 758
rect 1150 757 1158 758
rect 467 755 475 756
rect 325 751 333 752
rect 467 752 475 753
rect 1082 752 1090 753
rect 1172 752 1180 753
rect 1326 756 1334 757
rect 1416 756 1424 757
rect 1348 751 1356 752
rect 1438 751 1446 752
rect 1082 749 1090 750
rect 1172 749 1180 750
rect -159 730 -151 731
rect -69 730 -61 731
rect 107 729 115 730
rect 197 729 205 730
rect 1348 748 1356 749
rect 1438 748 1446 749
rect -159 727 -151 728
rect -69 727 -61 728
rect -137 722 -129 723
rect -47 722 -39 723
rect 107 726 115 727
rect 197 726 205 727
rect 129 721 137 722
rect 219 721 227 722
rect -137 719 -129 720
rect -47 719 -39 720
rect 129 718 137 719
rect 219 718 227 719
rect 359 713 367 714
rect 359 710 367 711
rect 381 705 389 706
rect -218 681 -210 682
rect 381 702 389 703
rect 48 680 56 681
rect -218 678 -210 679
rect -196 673 -188 674
rect 48 677 56 678
rect 70 672 78 673
rect -196 670 -188 671
rect 70 669 78 670
rect 1045 667 1046 675
rect 1048 667 1049 675
rect 784 657 785 665
rect 787 657 788 665
rect 819 637 827 638
rect 819 634 827 635
rect 1064 630 1072 631
rect 1154 630 1162 631
rect 841 629 849 630
rect 1330 629 1338 630
rect 1420 629 1428 630
rect 1064 627 1072 628
rect 1154 627 1162 628
rect 841 626 849 627
rect 1086 622 1094 623
rect 1176 622 1184 623
rect 1330 626 1338 627
rect 1420 626 1428 627
rect 1352 621 1360 622
rect 1442 621 1450 622
rect 1086 619 1094 620
rect 1176 619 1184 620
rect 314 600 322 601
rect 1352 618 1360 619
rect 1442 618 1450 619
rect 314 597 322 598
rect -163 588 -155 589
rect -73 588 -65 589
rect 103 587 111 588
rect 193 587 201 588
rect 336 592 344 593
rect 905 592 913 593
rect -163 585 -155 586
rect -73 585 -65 586
rect -141 580 -133 581
rect -51 580 -43 581
rect 103 584 111 585
rect 193 584 201 585
rect 336 589 344 590
rect 401 582 402 590
rect 404 582 405 590
rect 785 583 793 584
rect 905 589 913 590
rect 927 584 935 585
rect 125 579 133 580
rect 215 579 223 580
rect -141 577 -133 578
rect -51 577 -43 578
rect 785 580 793 581
rect 125 576 133 577
rect 215 576 223 577
rect 927 581 935 582
rect 1005 581 1013 582
rect 1271 580 1279 581
rect 1005 578 1013 579
rect 1027 573 1035 574
rect 1271 577 1279 578
rect 1293 572 1301 573
rect 1027 570 1035 571
rect 1293 569 1301 570
rect 819 542 827 543
rect 819 539 827 540
rect 841 534 849 535
rect 841 531 849 532
rect -178 495 -177 503
rect -175 495 -174 503
rect 324 493 325 501
rect 327 493 328 501
rect 1060 488 1068 489
rect 1150 488 1158 489
rect 1326 487 1334 488
rect 1416 487 1424 488
rect 1060 485 1068 486
rect 1150 485 1158 486
rect 1082 480 1090 481
rect 1172 480 1180 481
rect 1326 484 1334 485
rect 1416 484 1424 485
rect 359 473 367 474
rect 1348 479 1356 480
rect 1438 479 1446 480
rect 359 470 367 471
rect -159 458 -151 459
rect -69 458 -61 459
rect 1082 477 1090 478
rect 1172 477 1180 478
rect 381 465 389 466
rect 1348 476 1356 477
rect 1438 476 1446 477
rect 107 457 115 458
rect 197 457 205 458
rect -159 455 -151 456
rect -69 455 -61 456
rect -137 450 -129 451
rect -47 450 -39 451
rect 107 454 115 455
rect 197 454 205 455
rect 381 462 389 463
rect 129 449 137 450
rect 219 449 227 450
rect -137 447 -129 448
rect -47 447 -39 448
rect 129 446 137 447
rect 219 446 227 447
rect 445 428 453 429
rect -218 409 -210 410
rect 48 408 56 409
rect 325 419 333 420
rect 445 425 453 426
rect 467 420 475 421
rect 325 416 333 417
rect 467 417 475 418
rect -218 406 -210 407
rect -196 401 -188 402
rect 48 405 56 406
rect 70 400 78 401
rect -196 398 -188 399
rect 70 397 78 398
rect 1045 395 1046 403
rect 1048 395 1049 403
rect 359 378 367 379
rect 359 375 367 376
rect 381 370 389 371
rect 381 367 389 368
rect 1064 358 1072 359
rect 1154 358 1162 359
rect 1330 357 1338 358
rect 1420 357 1428 358
rect 1064 355 1072 356
rect 1154 355 1162 356
rect 1086 350 1094 351
rect 1176 350 1184 351
rect 1330 354 1338 355
rect 1420 354 1428 355
rect 1352 349 1360 350
rect 1442 349 1450 350
rect 1086 347 1094 348
rect 1176 347 1184 348
rect 1352 346 1360 347
rect 1442 346 1450 347
rect -163 316 -155 317
rect -73 316 -65 317
rect 103 315 111 316
rect 193 315 201 316
rect -163 313 -155 314
rect -73 313 -65 314
rect -141 308 -133 309
rect -51 308 -43 309
rect 103 312 111 313
rect 193 312 201 313
rect 1005 309 1013 310
rect 125 307 133 308
rect 215 307 223 308
rect 1271 308 1279 309
rect -141 305 -133 306
rect -51 305 -43 306
rect 1005 306 1013 307
rect 125 304 133 305
rect 215 304 223 305
rect 1027 301 1035 302
rect 1271 305 1279 306
rect 1293 300 1301 301
rect 1027 298 1035 299
rect 1293 297 1301 298
rect 314 265 322 266
rect 314 262 322 263
rect 336 257 344 258
rect 336 254 344 255
rect 401 247 402 255
rect 404 247 405 255
rect -178 223 -177 231
rect -175 223 -174 231
rect -159 186 -151 187
rect -69 186 -61 187
rect 107 185 115 186
rect 197 185 205 186
rect -159 183 -151 184
rect -69 183 -61 184
rect -137 178 -129 179
rect -47 178 -39 179
rect 107 182 115 183
rect 197 182 205 183
rect 129 177 137 178
rect 219 177 227 178
rect -137 175 -129 176
rect -47 175 -39 176
rect 129 174 137 175
rect 219 174 227 175
rect -218 137 -210 138
rect 48 136 56 137
rect -218 134 -210 135
rect -196 129 -188 130
rect 48 133 56 134
rect 70 128 78 129
rect -196 126 -188 127
rect 70 125 78 126
rect -163 44 -155 45
rect -73 44 -65 45
rect 103 43 111 44
rect 193 43 201 44
rect -163 41 -155 42
rect -73 41 -65 42
rect -141 36 -133 37
rect -51 36 -43 37
rect 103 40 111 41
rect 193 40 201 41
rect 125 35 133 36
rect 215 35 223 36
rect -141 33 -133 34
rect -51 33 -43 34
rect 125 32 133 33
rect 215 32 223 33
rect -178 -49 -177 -41
rect -175 -49 -174 -41
rect -159 -86 -151 -85
rect -69 -86 -61 -85
rect 107 -87 115 -86
rect 197 -87 205 -86
rect -159 -89 -151 -88
rect -69 -89 -61 -88
rect -137 -94 -129 -93
rect -47 -94 -39 -93
rect 107 -90 115 -89
rect 197 -90 205 -89
rect 129 -95 137 -94
rect 219 -95 227 -94
rect -137 -97 -129 -96
rect -47 -97 -39 -96
rect 129 -98 137 -97
rect 219 -98 227 -97
rect -218 -135 -210 -134
rect 48 -136 56 -135
rect -218 -138 -210 -137
rect -196 -143 -188 -142
rect 48 -139 56 -138
rect 70 -144 78 -143
rect -196 -146 -188 -145
rect 70 -147 78 -146
<< pdiffusion >>
rect -117 1966 -109 1967
rect -27 1966 -19 1967
rect 149 1965 157 1966
rect 239 1965 247 1966
rect -117 1963 -109 1964
rect -27 1963 -19 1964
rect 149 1962 157 1963
rect 239 1962 247 1963
rect -117 1914 -109 1915
rect -27 1914 -19 1915
rect 149 1913 157 1914
rect 239 1913 247 1914
rect -117 1911 -109 1912
rect -27 1911 -19 1912
rect 149 1910 157 1911
rect 239 1910 247 1911
rect -178 1875 -177 1883
rect -175 1875 -174 1883
rect -113 1836 -105 1837
rect -23 1836 -15 1837
rect 153 1835 161 1836
rect 243 1835 251 1836
rect -113 1833 -105 1834
rect -23 1833 -15 1834
rect 153 1832 161 1833
rect 243 1832 251 1833
rect -172 1787 -164 1788
rect -172 1784 -164 1785
rect -113 1784 -105 1785
rect 94 1786 102 1787
rect -23 1784 -15 1785
rect 94 1783 102 1784
rect 153 1783 161 1784
rect 243 1783 251 1784
rect -113 1781 -105 1782
rect -23 1781 -15 1782
rect 153 1780 161 1781
rect 243 1780 251 1781
rect -172 1735 -164 1736
rect 94 1734 102 1735
rect -172 1732 -164 1733
rect 94 1731 102 1732
rect -117 1694 -109 1695
rect -27 1694 -19 1695
rect 149 1693 157 1694
rect 239 1693 247 1694
rect -117 1691 -109 1692
rect -27 1691 -19 1692
rect 149 1690 157 1691
rect 239 1690 247 1691
rect -117 1642 -109 1643
rect -27 1642 -19 1643
rect 149 1641 157 1642
rect 239 1641 247 1642
rect -117 1639 -109 1640
rect -27 1639 -19 1640
rect 149 1638 157 1639
rect 239 1638 247 1639
rect -178 1603 -177 1611
rect -175 1603 -174 1611
rect 1106 1594 1114 1595
rect 1196 1594 1204 1595
rect 1372 1593 1380 1594
rect 1462 1593 1470 1594
rect 1106 1591 1114 1592
rect 1196 1591 1204 1592
rect 1372 1590 1380 1591
rect 1462 1590 1470 1591
rect -113 1564 -105 1565
rect -23 1564 -15 1565
rect 153 1563 161 1564
rect 243 1563 251 1564
rect -113 1561 -105 1562
rect -23 1561 -15 1562
rect 153 1560 161 1561
rect 243 1560 251 1561
rect 1106 1542 1114 1543
rect 1196 1542 1204 1543
rect 1372 1541 1380 1542
rect 1462 1541 1470 1542
rect 1106 1539 1114 1540
rect 1196 1539 1204 1540
rect 1372 1538 1380 1539
rect 1462 1538 1470 1539
rect -172 1515 -164 1516
rect -172 1512 -164 1513
rect -113 1512 -105 1513
rect 324 1518 325 1526
rect 327 1518 328 1526
rect 94 1514 102 1515
rect -23 1512 -15 1513
rect 94 1511 102 1512
rect 153 1511 161 1512
rect 243 1511 251 1512
rect -113 1509 -105 1510
rect -23 1509 -15 1510
rect 153 1508 161 1509
rect 243 1508 251 1509
rect 1045 1503 1046 1511
rect 1048 1503 1049 1511
rect 405 1496 413 1497
rect 405 1493 413 1494
rect -172 1463 -164 1464
rect 94 1462 102 1463
rect -172 1460 -164 1461
rect 94 1459 102 1460
rect 1110 1464 1118 1465
rect 1200 1464 1208 1465
rect 1376 1463 1384 1464
rect 1466 1463 1474 1464
rect 1110 1461 1118 1462
rect 1200 1461 1208 1462
rect 1376 1460 1384 1461
rect 1466 1460 1474 1461
rect 491 1451 499 1452
rect 405 1444 413 1445
rect 491 1448 499 1449
rect 405 1441 413 1442
rect -117 1422 -109 1423
rect -27 1422 -19 1423
rect 149 1421 157 1422
rect 345 1424 353 1425
rect 239 1421 247 1422
rect -117 1419 -109 1420
rect -27 1419 -19 1420
rect 149 1418 157 1419
rect 239 1418 247 1419
rect 345 1421 353 1422
rect 1051 1415 1059 1416
rect 1051 1412 1059 1413
rect 1110 1412 1118 1413
rect 1317 1414 1325 1415
rect 1200 1412 1208 1413
rect 1317 1411 1325 1412
rect 1376 1411 1384 1412
rect 1466 1411 1474 1412
rect 405 1401 413 1402
rect 1110 1409 1118 1410
rect 491 1399 499 1400
rect 405 1398 413 1399
rect 1200 1409 1208 1410
rect 1376 1408 1384 1409
rect 491 1396 499 1397
rect 1466 1408 1474 1409
rect 784 1376 785 1384
rect 787 1376 788 1384
rect -117 1370 -109 1371
rect -27 1370 -19 1371
rect 149 1369 157 1370
rect 239 1369 247 1370
rect -117 1367 -109 1368
rect -27 1367 -19 1368
rect 149 1366 157 1367
rect 239 1366 247 1367
rect 1051 1363 1059 1364
rect 1317 1362 1325 1363
rect 1051 1360 1059 1361
rect 865 1354 873 1355
rect 1317 1359 1325 1360
rect 405 1349 413 1350
rect 865 1351 873 1352
rect 405 1346 413 1347
rect -178 1331 -177 1339
rect -175 1331 -174 1339
rect 1106 1322 1114 1323
rect 1196 1322 1204 1323
rect 1372 1321 1380 1322
rect 1462 1321 1470 1322
rect 1106 1319 1114 1320
rect 1196 1319 1204 1320
rect 1372 1318 1380 1319
rect 1462 1318 1470 1319
rect 951 1309 959 1310
rect 865 1302 873 1303
rect 951 1306 959 1307
rect -113 1292 -105 1293
rect -23 1292 -15 1293
rect 865 1299 873 1300
rect 153 1291 161 1292
rect 243 1291 251 1292
rect -113 1289 -105 1290
rect -23 1289 -15 1290
rect 153 1288 161 1289
rect 243 1288 251 1289
rect 360 1288 368 1289
rect 360 1285 368 1286
rect 805 1282 813 1283
rect 401 1272 402 1280
rect 404 1272 405 1280
rect 805 1279 813 1280
rect 1106 1270 1114 1271
rect 1196 1270 1204 1271
rect 1372 1269 1380 1270
rect 1462 1269 1470 1270
rect 1106 1267 1114 1268
rect 865 1259 873 1260
rect 1196 1267 1204 1268
rect 1372 1266 1380 1267
rect 1462 1266 1470 1267
rect 951 1257 959 1258
rect 865 1256 873 1257
rect 951 1254 959 1255
rect -172 1243 -164 1244
rect -172 1240 -164 1241
rect -113 1240 -105 1241
rect 94 1242 102 1243
rect -23 1240 -15 1241
rect 94 1239 102 1240
rect 153 1239 161 1240
rect 243 1239 251 1240
rect -113 1237 -105 1238
rect -23 1237 -15 1238
rect 153 1236 161 1237
rect 243 1236 251 1237
rect 360 1236 368 1237
rect 360 1233 368 1234
rect 1045 1231 1046 1239
rect 1048 1231 1049 1239
rect 865 1207 873 1208
rect 865 1204 873 1205
rect -172 1191 -164 1192
rect 1110 1192 1118 1193
rect 1200 1192 1208 1193
rect 94 1190 102 1191
rect -172 1188 -164 1189
rect 94 1187 102 1188
rect 324 1183 325 1191
rect 327 1183 328 1191
rect 1376 1191 1384 1192
rect 1466 1191 1474 1192
rect 1110 1189 1118 1190
rect 1200 1189 1208 1190
rect 1376 1188 1384 1189
rect 1466 1188 1474 1189
rect 405 1161 413 1162
rect 405 1158 413 1159
rect -117 1150 -109 1151
rect -27 1150 -19 1151
rect 149 1149 157 1150
rect 239 1149 247 1150
rect -117 1147 -109 1148
rect -27 1147 -19 1148
rect 149 1146 157 1147
rect 239 1146 247 1147
rect 784 1143 785 1151
rect 787 1143 788 1151
rect 1051 1143 1059 1144
rect 1051 1140 1059 1141
rect 1110 1140 1118 1141
rect 1317 1142 1325 1143
rect 1200 1140 1208 1141
rect 1317 1139 1325 1140
rect 1376 1139 1384 1140
rect 1466 1139 1474 1140
rect 1110 1137 1118 1138
rect 1200 1137 1208 1138
rect 1376 1136 1384 1137
rect 1466 1136 1474 1137
rect 865 1121 873 1122
rect 491 1116 499 1117
rect 865 1118 873 1119
rect 405 1109 413 1110
rect 491 1113 499 1114
rect 405 1106 413 1107
rect -117 1098 -109 1099
rect -27 1098 -19 1099
rect 149 1097 157 1098
rect 239 1097 247 1098
rect -117 1095 -109 1096
rect -27 1095 -19 1096
rect 149 1094 157 1095
rect 239 1094 247 1095
rect 345 1089 353 1090
rect 345 1086 353 1087
rect 1051 1091 1059 1092
rect 1317 1090 1325 1091
rect 1051 1088 1059 1089
rect 1317 1087 1325 1088
rect 951 1076 959 1077
rect -178 1059 -177 1067
rect -175 1059 -174 1067
rect 865 1069 873 1070
rect 951 1073 959 1074
rect 405 1066 413 1067
rect 491 1064 499 1065
rect 405 1063 413 1064
rect 865 1066 873 1067
rect 491 1061 499 1062
rect 1106 1050 1114 1051
rect 1196 1050 1204 1051
rect 805 1049 813 1050
rect 1372 1049 1380 1050
rect 1462 1049 1470 1050
rect 805 1046 813 1047
rect 1106 1047 1114 1048
rect 1196 1047 1204 1048
rect 1372 1046 1380 1047
rect 1462 1046 1470 1047
rect -113 1020 -105 1021
rect -23 1020 -15 1021
rect 153 1019 161 1020
rect 546 1023 547 1031
rect 549 1023 550 1031
rect 584 1023 585 1031
rect 587 1023 588 1031
rect 622 1023 623 1031
rect 625 1023 626 1031
rect 660 1023 661 1031
rect 663 1023 664 1031
rect 729 1024 730 1032
rect 732 1024 733 1032
rect 865 1026 873 1027
rect 951 1024 959 1025
rect 243 1019 251 1020
rect -113 1017 -105 1018
rect -23 1017 -15 1018
rect 153 1016 161 1017
rect 243 1016 251 1017
rect 405 1014 413 1015
rect 405 1011 413 1012
rect 865 1023 873 1024
rect 951 1021 959 1022
rect 1106 998 1114 999
rect 1196 998 1204 999
rect 1372 997 1380 998
rect 1462 997 1470 998
rect 1106 995 1114 996
rect 1196 995 1204 996
rect 1372 994 1380 995
rect 1462 994 1470 995
rect -172 971 -164 972
rect -172 968 -164 969
rect -113 968 -105 969
rect 94 970 102 971
rect -23 968 -15 969
rect 94 967 102 968
rect 153 967 161 968
rect 243 967 251 968
rect -113 965 -105 966
rect -23 965 -15 966
rect 729 967 730 975
rect 732 967 733 975
rect 865 974 873 975
rect 865 971 873 972
rect 153 964 161 965
rect 243 964 251 965
rect 360 953 368 954
rect 1045 959 1046 967
rect 1048 959 1049 967
rect 360 950 368 951
rect 401 937 402 945
rect 404 937 405 945
rect -172 919 -164 920
rect 94 918 102 919
rect -172 916 -164 917
rect 94 915 102 916
rect 1110 920 1118 921
rect 1200 920 1208 921
rect 1376 919 1384 920
rect 1466 919 1474 920
rect 729 910 730 918
rect 732 910 733 918
rect 784 910 785 918
rect 787 910 788 918
rect 1110 917 1118 918
rect 1200 917 1208 918
rect 1376 916 1384 917
rect 1466 916 1474 917
rect 360 901 368 902
rect 360 898 368 899
rect -117 878 -109 879
rect -27 878 -19 879
rect 865 888 873 889
rect 149 877 157 878
rect 865 885 873 886
rect 239 877 247 878
rect -117 875 -109 876
rect -27 875 -19 876
rect 149 874 157 875
rect 239 874 247 875
rect 1051 871 1059 872
rect 1051 868 1059 869
rect 1110 868 1118 869
rect 1317 870 1325 871
rect 1200 868 1208 869
rect 1317 867 1325 868
rect 1376 867 1384 868
rect 1466 867 1474 868
rect 324 848 325 856
rect 327 848 328 856
rect 729 853 730 861
rect 732 853 733 861
rect 1110 865 1118 866
rect 1200 865 1208 866
rect 1376 864 1384 865
rect 1466 864 1474 865
rect 951 843 959 844
rect -117 826 -109 827
rect -27 826 -19 827
rect 149 825 157 826
rect 865 836 873 837
rect 951 840 959 841
rect 239 825 247 826
rect 865 833 873 834
rect 405 826 413 827
rect -117 823 -109 824
rect -27 823 -19 824
rect 405 823 413 824
rect 149 822 157 823
rect 239 822 247 823
rect 1051 819 1059 820
rect 1317 818 1325 819
rect 805 816 813 817
rect 805 813 813 814
rect 1051 816 1059 817
rect 1317 815 1325 816
rect -178 787 -177 795
rect -175 787 -174 795
rect 865 793 873 794
rect 951 791 959 792
rect 865 790 873 791
rect 951 788 959 789
rect 491 781 499 782
rect 405 774 413 775
rect 491 778 499 779
rect 1106 778 1114 779
rect 1196 778 1204 779
rect 1372 777 1380 778
rect 1462 777 1470 778
rect 1106 775 1114 776
rect 405 771 413 772
rect 1196 775 1204 776
rect 1372 774 1380 775
rect 1462 774 1470 775
rect -113 748 -105 749
rect -23 748 -15 749
rect 345 754 353 755
rect 153 747 161 748
rect 243 747 251 748
rect 345 751 353 752
rect -113 745 -105 746
rect -23 745 -15 746
rect 153 744 161 745
rect 243 744 251 745
rect 865 741 873 742
rect 865 738 873 739
rect 405 731 413 732
rect 491 729 499 730
rect 405 728 413 729
rect 491 726 499 727
rect 1106 726 1114 727
rect 1196 726 1204 727
rect 1372 725 1380 726
rect 1462 725 1470 726
rect 1106 723 1114 724
rect 1196 723 1204 724
rect 1372 722 1380 723
rect 1462 722 1470 723
rect -172 699 -164 700
rect -172 696 -164 697
rect -113 696 -105 697
rect 94 698 102 699
rect -23 696 -15 697
rect 94 695 102 696
rect 153 695 161 696
rect 243 695 251 696
rect -113 693 -105 694
rect -23 693 -15 694
rect 153 692 161 693
rect 243 692 251 693
rect 1045 687 1046 695
rect 1048 687 1049 695
rect 405 679 413 680
rect 784 677 785 685
rect 787 677 788 685
rect 405 676 413 677
rect 865 655 873 656
rect 865 652 873 653
rect -172 647 -164 648
rect 1110 648 1118 649
rect 1200 648 1208 649
rect 94 646 102 647
rect -172 644 -164 645
rect 94 643 102 644
rect 1376 647 1384 648
rect 1466 647 1474 648
rect 1110 645 1118 646
rect 1200 645 1208 646
rect 1376 644 1384 645
rect 1466 644 1474 645
rect 360 618 368 619
rect 360 615 368 616
rect -117 606 -109 607
rect -27 606 -19 607
rect 951 610 959 611
rect 149 605 157 606
rect 239 605 247 606
rect -117 603 -109 604
rect -27 603 -19 604
rect 149 602 157 603
rect 239 602 247 603
rect 401 602 402 610
rect 404 602 405 610
rect 865 603 873 604
rect 951 607 959 608
rect 865 600 873 601
rect 1051 599 1059 600
rect 1051 596 1059 597
rect 1110 596 1118 597
rect 1317 598 1325 599
rect 1200 596 1208 597
rect 1317 595 1325 596
rect 1376 595 1384 596
rect 1466 595 1474 596
rect 1110 593 1118 594
rect 805 583 813 584
rect 805 580 813 581
rect 1200 593 1208 594
rect 1376 592 1384 593
rect 1466 592 1474 593
rect 360 566 368 567
rect 360 563 368 564
rect -117 554 -109 555
rect -27 554 -19 555
rect 149 553 157 554
rect 865 560 873 561
rect 951 558 959 559
rect 865 557 873 558
rect 239 553 247 554
rect -117 551 -109 552
rect -27 551 -19 552
rect 951 555 959 556
rect 149 550 157 551
rect 239 550 247 551
rect 1051 547 1059 548
rect 1317 546 1325 547
rect 1051 544 1059 545
rect 1317 543 1325 544
rect -178 515 -177 523
rect -175 515 -174 523
rect 324 513 325 521
rect 327 513 328 521
rect 865 508 873 509
rect 1106 506 1114 507
rect 1196 506 1204 507
rect 865 505 873 506
rect 1372 505 1380 506
rect 1462 505 1470 506
rect 1106 503 1114 504
rect 1196 503 1204 504
rect 1372 502 1380 503
rect 1462 502 1470 503
rect 405 491 413 492
rect 405 488 413 489
rect -113 476 -105 477
rect -23 476 -15 477
rect 153 475 161 476
rect 243 475 251 476
rect -113 473 -105 474
rect -23 473 -15 474
rect 153 472 161 473
rect 243 472 251 473
rect 1106 454 1114 455
rect 1196 454 1204 455
rect 1372 453 1380 454
rect 1462 453 1470 454
rect 1106 451 1114 452
rect 491 446 499 447
rect 1196 451 1204 452
rect 1372 450 1380 451
rect 405 439 413 440
rect 491 443 499 444
rect 1462 450 1470 451
rect 405 436 413 437
rect -172 427 -164 428
rect -172 424 -164 425
rect -113 424 -105 425
rect 94 426 102 427
rect -23 424 -15 425
rect 94 423 102 424
rect 153 423 161 424
rect 243 423 251 424
rect -113 421 -105 422
rect -23 421 -15 422
rect 153 420 161 421
rect 243 420 251 421
rect 345 419 353 420
rect 345 416 353 417
rect 1045 415 1046 423
rect 1048 415 1049 423
rect 405 396 413 397
rect 491 394 499 395
rect 405 393 413 394
rect 491 391 499 392
rect -172 375 -164 376
rect 1110 376 1118 377
rect 1200 376 1208 377
rect 94 374 102 375
rect -172 372 -164 373
rect 94 371 102 372
rect 1376 375 1384 376
rect 1466 375 1474 376
rect 1110 373 1118 374
rect 1200 373 1208 374
rect 1376 372 1384 373
rect 1466 372 1474 373
rect 405 344 413 345
rect -117 334 -109 335
rect -27 334 -19 335
rect 405 341 413 342
rect 149 333 157 334
rect 239 333 247 334
rect -117 331 -109 332
rect -27 331 -19 332
rect 149 330 157 331
rect 239 330 247 331
rect 1051 327 1059 328
rect 1051 324 1059 325
rect 1110 324 1118 325
rect 1317 326 1325 327
rect 1200 324 1208 325
rect 1317 323 1325 324
rect 1376 323 1384 324
rect 1466 323 1474 324
rect 1110 321 1118 322
rect 1200 321 1208 322
rect 1376 320 1384 321
rect 1466 320 1474 321
rect -117 282 -109 283
rect -27 282 -19 283
rect 149 281 157 282
rect 360 283 368 284
rect 239 281 247 282
rect -117 279 -109 280
rect -27 279 -19 280
rect 360 280 368 281
rect 149 278 157 279
rect 239 278 247 279
rect 1051 275 1059 276
rect 401 267 402 275
rect 404 267 405 275
rect 1317 274 1325 275
rect 1051 272 1059 273
rect 1317 271 1325 272
rect -178 243 -177 251
rect -175 243 -174 251
rect 360 231 368 232
rect 360 228 368 229
rect -113 204 -105 205
rect -23 204 -15 205
rect 153 203 161 204
rect 243 203 251 204
rect -113 201 -105 202
rect -23 201 -15 202
rect 153 200 161 201
rect 243 200 251 201
rect -172 155 -164 156
rect -172 152 -164 153
rect -113 152 -105 153
rect 94 154 102 155
rect -23 152 -15 153
rect 94 151 102 152
rect 153 151 161 152
rect 243 151 251 152
rect -113 149 -105 150
rect -23 149 -15 150
rect 153 148 161 149
rect 243 148 251 149
rect -172 103 -164 104
rect 94 102 102 103
rect -172 100 -164 101
rect 94 99 102 100
rect -117 62 -109 63
rect -27 62 -19 63
rect 149 61 157 62
rect 239 61 247 62
rect -117 59 -109 60
rect -27 59 -19 60
rect 149 58 157 59
rect 239 58 247 59
rect -117 10 -109 11
rect -27 10 -19 11
rect 149 9 157 10
rect 239 9 247 10
rect -117 7 -109 8
rect -27 7 -19 8
rect 149 6 157 7
rect 239 6 247 7
rect -178 -29 -177 -21
rect -175 -29 -174 -21
rect -113 -68 -105 -67
rect -23 -68 -15 -67
rect 153 -69 161 -68
rect 243 -69 251 -68
rect -113 -71 -105 -70
rect -23 -71 -15 -70
rect 153 -72 161 -71
rect 243 -72 251 -71
rect -172 -117 -164 -116
rect -172 -120 -164 -119
rect -113 -120 -105 -119
rect 94 -118 102 -117
rect -23 -120 -15 -119
rect 94 -121 102 -120
rect 153 -121 161 -120
rect 243 -121 251 -120
rect -113 -123 -105 -122
rect -23 -123 -15 -122
rect 153 -124 161 -123
rect 243 -124 251 -123
rect -172 -169 -164 -168
rect 94 -170 102 -169
rect -172 -172 -164 -171
rect 94 -173 102 -172
<< ndcontact >>
rect -163 1949 -155 1953
rect -73 1949 -65 1953
rect 103 1948 111 1952
rect 193 1948 201 1952
rect -163 1941 -155 1945
rect -141 1941 -133 1945
rect -73 1941 -65 1945
rect -51 1941 -43 1945
rect 103 1940 111 1944
rect 125 1940 133 1944
rect 193 1940 201 1944
rect 215 1940 223 1944
rect -141 1933 -133 1937
rect -51 1933 -43 1937
rect 125 1932 133 1936
rect 215 1932 223 1936
rect -182 1855 -178 1863
rect -174 1855 -170 1863
rect -159 1819 -151 1823
rect -69 1819 -61 1823
rect 107 1818 115 1822
rect 197 1818 205 1822
rect -159 1811 -151 1815
rect -137 1811 -129 1815
rect -69 1811 -61 1815
rect -47 1811 -39 1815
rect 107 1810 115 1814
rect 129 1810 137 1814
rect 197 1810 205 1814
rect 219 1810 227 1814
rect -137 1803 -129 1807
rect -47 1803 -39 1807
rect 129 1802 137 1806
rect 219 1802 227 1806
rect -218 1770 -210 1774
rect 48 1769 56 1773
rect -218 1762 -210 1766
rect -196 1762 -188 1766
rect 48 1761 56 1765
rect 70 1761 78 1765
rect -196 1754 -188 1758
rect 70 1753 78 1757
rect -163 1677 -155 1681
rect -73 1677 -65 1681
rect 103 1676 111 1680
rect 193 1676 201 1680
rect -163 1669 -155 1673
rect -141 1669 -133 1673
rect -73 1669 -65 1673
rect -51 1669 -43 1673
rect 103 1668 111 1672
rect 125 1668 133 1672
rect 193 1668 201 1672
rect 215 1668 223 1672
rect -141 1661 -133 1665
rect -51 1661 -43 1665
rect 125 1660 133 1664
rect 215 1660 223 1664
rect -182 1583 -178 1591
rect -174 1583 -170 1591
rect 1060 1577 1068 1581
rect 1150 1577 1158 1581
rect 1326 1576 1334 1580
rect 1416 1576 1424 1580
rect 1060 1569 1068 1573
rect 1082 1569 1090 1573
rect 1150 1569 1158 1573
rect 1172 1569 1180 1573
rect 1326 1568 1334 1572
rect 1348 1568 1356 1572
rect 1416 1568 1424 1572
rect 1438 1568 1446 1572
rect 1082 1561 1090 1565
rect 1172 1561 1180 1565
rect -159 1547 -151 1551
rect -69 1547 -61 1551
rect 1348 1560 1356 1564
rect 1438 1560 1446 1564
rect 107 1546 115 1550
rect 197 1546 205 1550
rect -159 1539 -151 1543
rect -137 1539 -129 1543
rect -69 1539 -61 1543
rect -47 1539 -39 1543
rect 107 1538 115 1542
rect 129 1538 137 1542
rect 197 1538 205 1542
rect 219 1538 227 1542
rect -137 1531 -129 1535
rect -47 1531 -39 1535
rect 129 1530 137 1534
rect 219 1530 227 1534
rect -218 1498 -210 1502
rect 48 1497 56 1501
rect 320 1498 324 1506
rect 328 1498 332 1506
rect -218 1490 -210 1494
rect -196 1490 -188 1494
rect 48 1489 56 1493
rect 70 1489 78 1493
rect -196 1482 -188 1486
rect 70 1481 78 1485
rect 359 1479 367 1483
rect 1041 1483 1045 1491
rect 1049 1483 1053 1491
rect 359 1471 367 1475
rect 381 1471 389 1475
rect 381 1463 389 1467
rect 1064 1447 1072 1451
rect 1154 1447 1162 1451
rect 1330 1446 1338 1450
rect 1420 1446 1428 1450
rect 1064 1439 1072 1443
rect 1086 1439 1094 1443
rect 1154 1439 1162 1443
rect 1176 1439 1184 1443
rect 445 1434 453 1438
rect 1330 1438 1338 1442
rect 1352 1438 1360 1442
rect 1420 1438 1428 1442
rect 1442 1438 1450 1442
rect 325 1425 333 1429
rect 445 1426 453 1430
rect 467 1426 475 1430
rect 1086 1431 1094 1435
rect 1176 1431 1184 1435
rect 1352 1430 1360 1434
rect 1442 1430 1450 1434
rect 325 1417 333 1421
rect 467 1418 475 1422
rect -163 1405 -155 1409
rect -73 1405 -65 1409
rect 103 1404 111 1408
rect 193 1404 201 1408
rect -163 1397 -155 1401
rect -141 1397 -133 1401
rect -73 1397 -65 1401
rect -51 1397 -43 1401
rect 103 1396 111 1400
rect 125 1396 133 1400
rect 193 1396 201 1400
rect 215 1396 223 1400
rect -141 1389 -133 1393
rect 1005 1398 1013 1402
rect 1271 1397 1279 1401
rect -51 1389 -43 1393
rect 125 1388 133 1392
rect 215 1388 223 1392
rect 1005 1390 1013 1394
rect 1027 1390 1035 1394
rect 1271 1389 1279 1393
rect 1293 1389 1301 1393
rect 359 1384 367 1388
rect 359 1376 367 1380
rect 381 1376 389 1380
rect 1027 1382 1035 1386
rect 381 1368 389 1372
rect 1293 1381 1301 1385
rect 780 1356 784 1364
rect 788 1356 792 1364
rect 819 1337 827 1341
rect 819 1329 827 1333
rect 841 1329 849 1333
rect -182 1311 -178 1319
rect -174 1311 -170 1319
rect 841 1321 849 1325
rect 1060 1305 1068 1309
rect 1150 1305 1158 1309
rect 1326 1304 1334 1308
rect 1416 1304 1424 1308
rect 1060 1297 1068 1301
rect 1082 1297 1090 1301
rect 1150 1297 1158 1301
rect 1172 1297 1180 1301
rect 905 1292 913 1296
rect 1326 1296 1334 1300
rect 1348 1296 1356 1300
rect 1416 1296 1424 1300
rect 1438 1296 1446 1300
rect -159 1275 -151 1279
rect -69 1275 -61 1279
rect 785 1283 793 1287
rect 905 1284 913 1288
rect 927 1284 935 1288
rect 1082 1289 1090 1293
rect 1172 1289 1180 1293
rect 1348 1288 1356 1292
rect 1438 1288 1446 1292
rect 107 1274 115 1278
rect 197 1274 205 1278
rect 314 1271 322 1275
rect -159 1267 -151 1271
rect -137 1267 -129 1271
rect -69 1267 -61 1271
rect -47 1267 -39 1271
rect 785 1275 793 1279
rect 927 1276 935 1280
rect 107 1266 115 1270
rect 129 1266 137 1270
rect 197 1266 205 1270
rect 219 1266 227 1270
rect -137 1259 -129 1263
rect 314 1263 322 1267
rect 336 1263 344 1267
rect -47 1259 -39 1263
rect 129 1258 137 1262
rect 219 1258 227 1262
rect 336 1255 344 1259
rect 397 1252 401 1260
rect 405 1252 409 1260
rect 819 1242 827 1246
rect -218 1226 -210 1230
rect 48 1225 56 1229
rect 819 1234 827 1238
rect 841 1234 849 1238
rect 841 1226 849 1230
rect -218 1218 -210 1222
rect -196 1218 -188 1222
rect 48 1217 56 1221
rect 70 1217 78 1221
rect -196 1210 -188 1214
rect 70 1209 78 1213
rect 1041 1211 1045 1219
rect 1049 1211 1053 1219
rect 1064 1175 1072 1179
rect 1154 1175 1162 1179
rect 1330 1174 1338 1178
rect 1420 1174 1428 1178
rect 320 1163 324 1171
rect 328 1163 332 1171
rect 1064 1167 1072 1171
rect 1086 1167 1094 1171
rect 1154 1167 1162 1171
rect 1176 1167 1184 1171
rect 1330 1166 1338 1170
rect 1352 1166 1360 1170
rect 1420 1166 1428 1170
rect 1442 1166 1450 1170
rect 1086 1159 1094 1163
rect 1176 1159 1184 1163
rect 1352 1158 1360 1162
rect 1442 1158 1450 1162
rect 359 1144 367 1148
rect -163 1133 -155 1137
rect -73 1133 -65 1137
rect 103 1132 111 1136
rect 193 1132 201 1136
rect 359 1136 367 1140
rect 381 1136 389 1140
rect -163 1125 -155 1129
rect -141 1125 -133 1129
rect -73 1125 -65 1129
rect -51 1125 -43 1129
rect 103 1124 111 1128
rect 125 1124 133 1128
rect 193 1124 201 1128
rect 215 1124 223 1128
rect 381 1128 389 1132
rect -141 1117 -133 1121
rect -51 1117 -43 1121
rect 125 1116 133 1120
rect 780 1123 784 1131
rect 788 1123 792 1131
rect 1005 1126 1013 1130
rect 215 1116 223 1120
rect 1271 1125 1279 1129
rect 1005 1118 1013 1122
rect 1027 1118 1035 1122
rect 1271 1117 1279 1121
rect 1293 1117 1301 1121
rect 819 1104 827 1108
rect 445 1099 453 1103
rect 1027 1110 1035 1114
rect 1293 1109 1301 1113
rect 325 1090 333 1094
rect 819 1096 827 1100
rect 841 1096 849 1100
rect 445 1091 453 1095
rect 467 1091 475 1095
rect 325 1082 333 1086
rect 467 1083 475 1087
rect 841 1088 849 1092
rect 905 1059 913 1063
rect 359 1049 367 1053
rect 785 1050 793 1054
rect 905 1051 913 1055
rect 927 1051 935 1055
rect -182 1039 -178 1047
rect -174 1039 -170 1047
rect 359 1041 367 1045
rect 381 1041 389 1045
rect 785 1042 793 1046
rect 927 1043 935 1047
rect 381 1033 389 1037
rect 1060 1033 1068 1037
rect 1150 1033 1158 1037
rect 1326 1032 1334 1036
rect 1416 1032 1424 1036
rect 1060 1025 1068 1029
rect 1082 1025 1090 1029
rect 1150 1025 1158 1029
rect 1172 1025 1180 1029
rect 1326 1024 1334 1028
rect 1348 1024 1356 1028
rect 1416 1024 1424 1028
rect 1438 1024 1446 1028
rect -159 1003 -151 1007
rect -69 1003 -61 1007
rect 107 1002 115 1006
rect 197 1002 205 1006
rect 725 1004 729 1012
rect 733 1004 737 1012
rect 819 1009 827 1013
rect 1082 1017 1090 1021
rect 1172 1017 1180 1021
rect 1348 1016 1356 1020
rect 1438 1016 1446 1020
rect 819 1001 827 1005
rect 841 1001 849 1005
rect -159 995 -151 999
rect -137 995 -129 999
rect -69 995 -61 999
rect -47 995 -39 999
rect 107 994 115 998
rect 129 994 137 998
rect 197 994 205 998
rect 219 994 227 998
rect -137 987 -129 991
rect -47 987 -39 991
rect 129 986 137 990
rect 219 986 227 990
rect 656 983 660 991
rect 664 983 668 991
rect 686 984 690 992
rect 694 984 698 992
rect 841 993 849 997
rect -218 954 -210 958
rect 48 953 56 957
rect 648 953 652 961
rect 656 953 660 961
rect -218 946 -210 950
rect -196 946 -188 950
rect 48 945 56 949
rect 70 945 78 949
rect -196 938 -188 942
rect 70 937 78 941
rect 314 936 322 940
rect 618 942 622 950
rect 626 942 630 950
rect 725 947 729 955
rect 733 947 737 955
rect 1041 939 1045 947
rect 1049 939 1053 947
rect 314 928 322 932
rect 336 928 344 932
rect 336 920 344 924
rect 397 917 401 925
rect 405 917 409 925
rect 610 912 614 920
rect 618 912 622 920
rect 580 901 584 909
rect 588 901 592 909
rect 1064 903 1072 907
rect 1154 903 1162 907
rect 1330 902 1338 906
rect 1420 902 1428 906
rect 725 890 729 898
rect 733 890 737 898
rect 780 890 784 898
rect 788 890 792 898
rect 1064 895 1072 899
rect 1086 895 1094 899
rect 1154 895 1162 899
rect 1176 895 1184 899
rect 1330 894 1338 898
rect 1352 894 1360 898
rect 1420 894 1428 898
rect 1442 894 1450 898
rect 1086 887 1094 891
rect 1176 887 1184 891
rect -163 861 -155 865
rect -73 861 -65 865
rect 572 871 576 879
rect 580 871 584 879
rect 1352 886 1360 890
rect 1442 886 1450 890
rect 819 871 827 875
rect 103 860 111 864
rect 193 860 201 864
rect 542 860 546 868
rect 550 860 554 868
rect 819 863 827 867
rect 841 863 849 867
rect -163 853 -155 857
rect -141 853 -133 857
rect -73 853 -65 857
rect -51 853 -43 857
rect 103 852 111 856
rect 125 852 133 856
rect 193 852 201 856
rect 215 852 223 856
rect -141 845 -133 849
rect -51 845 -43 849
rect 125 844 133 848
rect 215 844 223 848
rect 841 855 849 859
rect 1005 854 1013 858
rect 1271 853 1279 857
rect 1005 846 1013 850
rect 1027 846 1035 850
rect 1271 845 1279 849
rect 1293 845 1301 849
rect 320 828 324 836
rect 328 828 332 836
rect 534 831 538 839
rect 542 831 546 839
rect 725 833 729 841
rect 733 833 737 841
rect 1027 838 1035 842
rect 905 826 913 830
rect 1293 837 1301 841
rect 785 817 793 821
rect 905 818 913 822
rect 927 818 935 822
rect 359 809 367 813
rect 359 801 367 805
rect 381 801 389 805
rect 526 802 530 810
rect 534 802 538 810
rect 785 809 793 813
rect 927 810 935 814
rect 381 793 389 797
rect -182 767 -178 775
rect -174 767 -170 775
rect 819 776 827 780
rect 445 764 453 768
rect 819 768 827 772
rect 841 768 849 772
rect 325 755 333 759
rect 445 756 453 760
rect 467 756 475 760
rect 841 760 849 764
rect 1060 761 1068 765
rect 1150 761 1158 765
rect 1326 760 1334 764
rect 1416 760 1424 764
rect 325 747 333 751
rect 1060 753 1068 757
rect 1082 753 1090 757
rect 1150 753 1158 757
rect 1172 753 1180 757
rect 1326 752 1334 756
rect 1348 752 1356 756
rect 1416 752 1424 756
rect 1438 752 1446 756
rect 467 748 475 752
rect 1082 745 1090 749
rect 1172 745 1180 749
rect -159 731 -151 735
rect -69 731 -61 735
rect 107 730 115 734
rect 197 730 205 734
rect 1348 744 1356 748
rect 1438 744 1446 748
rect -159 723 -151 727
rect -137 723 -129 727
rect -69 723 -61 727
rect -47 723 -39 727
rect 107 722 115 726
rect 129 722 137 726
rect 197 722 205 726
rect 219 722 227 726
rect -137 715 -129 719
rect -47 715 -39 719
rect 129 714 137 718
rect 219 714 227 718
rect 359 714 367 718
rect 359 706 367 710
rect 381 706 389 710
rect -218 682 -210 686
rect 381 698 389 702
rect 48 681 56 685
rect -218 674 -210 678
rect -196 674 -188 678
rect 48 673 56 677
rect 70 673 78 677
rect -196 666 -188 670
rect 70 665 78 669
rect 1041 667 1045 675
rect 1049 667 1053 675
rect 780 657 784 665
rect 788 657 792 665
rect 819 638 827 642
rect 819 630 827 634
rect 841 630 849 634
rect 1064 631 1072 635
rect 1154 631 1162 635
rect 1330 630 1338 634
rect 1420 630 1428 634
rect 841 622 849 626
rect 1064 623 1072 627
rect 1086 623 1094 627
rect 1154 623 1162 627
rect 1176 623 1184 627
rect 1330 622 1338 626
rect 1352 622 1360 626
rect 1420 622 1428 626
rect 1442 622 1450 626
rect 1086 615 1094 619
rect 1176 615 1184 619
rect 314 601 322 605
rect 1352 614 1360 618
rect 1442 614 1450 618
rect -163 589 -155 593
rect -73 589 -65 593
rect 314 593 322 597
rect 336 593 344 597
rect 103 588 111 592
rect 193 588 201 592
rect 905 593 913 597
rect -163 581 -155 585
rect -141 581 -133 585
rect -73 581 -65 585
rect -51 581 -43 585
rect 103 580 111 584
rect 125 580 133 584
rect 193 580 201 584
rect 215 580 223 584
rect 336 585 344 589
rect 397 582 401 590
rect 405 582 409 590
rect 785 584 793 588
rect 905 585 913 589
rect 927 585 935 589
rect -141 573 -133 577
rect 1005 582 1013 586
rect -51 573 -43 577
rect 125 572 133 576
rect 785 576 793 580
rect 215 572 223 576
rect 1271 581 1279 585
rect 927 577 935 581
rect 1005 574 1013 578
rect 1027 574 1035 578
rect 1271 573 1279 577
rect 1293 573 1301 577
rect 1027 566 1035 570
rect 1293 565 1301 569
rect 819 543 827 547
rect 819 535 827 539
rect 841 535 849 539
rect 841 527 849 531
rect -182 495 -178 503
rect -174 495 -170 503
rect 320 493 324 501
rect 328 493 332 501
rect 1060 489 1068 493
rect 1150 489 1158 493
rect 1326 488 1334 492
rect 1416 488 1424 492
rect 1060 481 1068 485
rect 1082 481 1090 485
rect 1150 481 1158 485
rect 1172 481 1180 485
rect 1326 480 1334 484
rect 1348 480 1356 484
rect 1416 480 1424 484
rect 1438 480 1446 484
rect 359 474 367 478
rect -159 459 -151 463
rect -69 459 -61 463
rect 359 466 367 470
rect 381 466 389 470
rect 1082 473 1090 477
rect 1172 473 1180 477
rect 1348 472 1356 476
rect 1438 472 1446 476
rect 107 458 115 462
rect 197 458 205 462
rect -159 451 -151 455
rect -137 451 -129 455
rect -69 451 -61 455
rect -47 451 -39 455
rect 381 458 389 462
rect 107 450 115 454
rect 129 450 137 454
rect 197 450 205 454
rect 219 450 227 454
rect -137 443 -129 447
rect -47 443 -39 447
rect 129 442 137 446
rect 219 442 227 446
rect 445 429 453 433
rect -218 410 -210 414
rect 48 409 56 413
rect 325 420 333 424
rect 445 421 453 425
rect 467 421 475 425
rect 325 412 333 416
rect 467 413 475 417
rect -218 402 -210 406
rect -196 402 -188 406
rect 48 401 56 405
rect 70 401 78 405
rect -196 394 -188 398
rect 70 393 78 397
rect 1041 395 1045 403
rect 1049 395 1053 403
rect 359 379 367 383
rect 359 371 367 375
rect 381 371 389 375
rect 381 363 389 367
rect 1064 359 1072 363
rect 1154 359 1162 363
rect 1330 358 1338 362
rect 1420 358 1428 362
rect 1064 351 1072 355
rect 1086 351 1094 355
rect 1154 351 1162 355
rect 1176 351 1184 355
rect 1330 350 1338 354
rect 1352 350 1360 354
rect 1420 350 1428 354
rect 1442 350 1450 354
rect 1086 343 1094 347
rect 1176 343 1184 347
rect 1352 342 1360 346
rect 1442 342 1450 346
rect -163 317 -155 321
rect -73 317 -65 321
rect 103 316 111 320
rect 193 316 201 320
rect -163 309 -155 313
rect -141 309 -133 313
rect -73 309 -65 313
rect -51 309 -43 313
rect 103 308 111 312
rect 125 308 133 312
rect 193 308 201 312
rect 215 308 223 312
rect 1005 310 1013 314
rect 1271 309 1279 313
rect -141 301 -133 305
rect -51 301 -43 305
rect 125 300 133 304
rect 215 300 223 304
rect 1005 302 1013 306
rect 1027 302 1035 306
rect 1271 301 1279 305
rect 1293 301 1301 305
rect 1027 294 1035 298
rect 1293 293 1301 297
rect 314 266 322 270
rect 314 258 322 262
rect 336 258 344 262
rect 336 250 344 254
rect 397 247 401 255
rect 405 247 409 255
rect -182 223 -178 231
rect -174 223 -170 231
rect -159 187 -151 191
rect -69 187 -61 191
rect 107 186 115 190
rect 197 186 205 190
rect -159 179 -151 183
rect -137 179 -129 183
rect -69 179 -61 183
rect -47 179 -39 183
rect 107 178 115 182
rect 129 178 137 182
rect 197 178 205 182
rect 219 178 227 182
rect -137 171 -129 175
rect -47 171 -39 175
rect 129 170 137 174
rect 219 170 227 174
rect -218 138 -210 142
rect 48 137 56 141
rect -218 130 -210 134
rect -196 130 -188 134
rect 48 129 56 133
rect 70 129 78 133
rect -196 122 -188 126
rect 70 121 78 125
rect -163 45 -155 49
rect -73 45 -65 49
rect 103 44 111 48
rect 193 44 201 48
rect -163 37 -155 41
rect -141 37 -133 41
rect -73 37 -65 41
rect -51 37 -43 41
rect 103 36 111 40
rect 125 36 133 40
rect 193 36 201 40
rect 215 36 223 40
rect -141 29 -133 33
rect -51 29 -43 33
rect 125 28 133 32
rect 215 28 223 32
rect -182 -49 -178 -41
rect -174 -49 -170 -41
rect -159 -85 -151 -81
rect -69 -85 -61 -81
rect 107 -86 115 -82
rect 197 -86 205 -82
rect -159 -93 -151 -89
rect -137 -93 -129 -89
rect -69 -93 -61 -89
rect -47 -93 -39 -89
rect 107 -94 115 -90
rect 129 -94 137 -90
rect 197 -94 205 -90
rect 219 -94 227 -90
rect -137 -101 -129 -97
rect -47 -101 -39 -97
rect 129 -102 137 -98
rect 219 -102 227 -98
rect -218 -134 -210 -130
rect 48 -135 56 -131
rect -218 -142 -210 -138
rect -196 -142 -188 -138
rect 48 -143 56 -139
rect 70 -143 78 -139
rect -196 -150 -188 -146
rect 70 -151 78 -147
<< pdcontact >>
rect -117 1967 -109 1971
rect -27 1967 -19 1971
rect 149 1966 157 1970
rect 239 1966 247 1970
rect -117 1959 -109 1963
rect -27 1959 -19 1963
rect 149 1958 157 1962
rect 239 1958 247 1962
rect -117 1915 -109 1919
rect -27 1915 -19 1919
rect 149 1914 157 1918
rect 239 1914 247 1918
rect -117 1907 -109 1911
rect -27 1907 -19 1911
rect 149 1906 157 1910
rect 239 1906 247 1910
rect -182 1875 -178 1883
rect -174 1875 -170 1883
rect -113 1837 -105 1841
rect -23 1837 -15 1841
rect 153 1836 161 1840
rect 243 1836 251 1840
rect -113 1829 -105 1833
rect -23 1829 -15 1833
rect 153 1828 161 1832
rect 243 1828 251 1832
rect -172 1788 -164 1792
rect -113 1785 -105 1789
rect -23 1785 -15 1789
rect 94 1787 102 1791
rect 153 1784 161 1788
rect -172 1780 -164 1784
rect 243 1784 251 1788
rect -113 1777 -105 1781
rect -23 1777 -15 1781
rect 94 1779 102 1783
rect 153 1776 161 1780
rect 243 1776 251 1780
rect -172 1736 -164 1740
rect 94 1735 102 1739
rect -172 1728 -164 1732
rect 94 1727 102 1731
rect -117 1695 -109 1699
rect -27 1695 -19 1699
rect 149 1694 157 1698
rect 239 1694 247 1698
rect -117 1687 -109 1691
rect -27 1687 -19 1691
rect 149 1686 157 1690
rect 239 1686 247 1690
rect -117 1643 -109 1647
rect -27 1643 -19 1647
rect 149 1642 157 1646
rect 239 1642 247 1646
rect -117 1635 -109 1639
rect -27 1635 -19 1639
rect 149 1634 157 1638
rect 239 1634 247 1638
rect -182 1603 -178 1611
rect -174 1603 -170 1611
rect 1106 1595 1114 1599
rect 1196 1595 1204 1599
rect 1372 1594 1380 1598
rect 1462 1594 1470 1598
rect 1106 1587 1114 1591
rect 1196 1587 1204 1591
rect 1372 1586 1380 1590
rect 1462 1586 1470 1590
rect -113 1565 -105 1569
rect -23 1565 -15 1569
rect 153 1564 161 1568
rect 243 1564 251 1568
rect -113 1557 -105 1561
rect -23 1557 -15 1561
rect 153 1556 161 1560
rect 243 1556 251 1560
rect 1106 1543 1114 1547
rect 1196 1543 1204 1547
rect 1372 1542 1380 1546
rect 1462 1542 1470 1546
rect 1106 1535 1114 1539
rect 1196 1535 1204 1539
rect 1372 1534 1380 1538
rect 1462 1534 1470 1538
rect -172 1516 -164 1520
rect -113 1513 -105 1517
rect -23 1513 -15 1517
rect 94 1515 102 1519
rect 320 1518 324 1526
rect 328 1518 332 1526
rect 153 1512 161 1516
rect -172 1508 -164 1512
rect 243 1512 251 1516
rect -113 1505 -105 1509
rect -23 1505 -15 1509
rect 94 1507 102 1511
rect 153 1504 161 1508
rect 243 1504 251 1508
rect 1041 1503 1045 1511
rect 1049 1503 1053 1511
rect 405 1497 413 1501
rect 405 1489 413 1493
rect -172 1464 -164 1468
rect 94 1463 102 1467
rect -172 1456 -164 1460
rect 1110 1465 1118 1469
rect 1200 1465 1208 1469
rect 1376 1464 1384 1468
rect 1466 1464 1474 1468
rect 94 1455 102 1459
rect 1110 1457 1118 1461
rect 1200 1457 1208 1461
rect 1376 1456 1384 1460
rect 1466 1456 1474 1460
rect 491 1452 499 1456
rect 405 1445 413 1449
rect 491 1444 499 1448
rect 405 1437 413 1441
rect -117 1423 -109 1427
rect -27 1423 -19 1427
rect 149 1422 157 1426
rect 239 1422 247 1426
rect 345 1425 353 1429
rect -117 1415 -109 1419
rect -27 1415 -19 1419
rect 149 1414 157 1418
rect 239 1414 247 1418
rect 345 1417 353 1421
rect 1051 1416 1059 1420
rect 1110 1413 1118 1417
rect 1200 1413 1208 1417
rect 1317 1415 1325 1419
rect 1376 1412 1384 1416
rect 1051 1408 1059 1412
rect 1466 1412 1474 1416
rect 405 1402 413 1406
rect 491 1400 499 1404
rect 405 1394 413 1398
rect 1110 1405 1118 1409
rect 1200 1405 1208 1409
rect 1317 1407 1325 1411
rect 491 1392 499 1396
rect 1376 1404 1384 1408
rect 1466 1404 1474 1408
rect 780 1376 784 1384
rect 788 1376 792 1384
rect -117 1371 -109 1375
rect -27 1371 -19 1375
rect 149 1370 157 1374
rect 239 1370 247 1374
rect -117 1363 -109 1367
rect -27 1363 -19 1367
rect 149 1362 157 1366
rect 239 1362 247 1366
rect 1051 1364 1059 1368
rect 1317 1363 1325 1367
rect 405 1350 413 1354
rect 865 1355 873 1359
rect 1051 1356 1059 1360
rect 1317 1355 1325 1359
rect 865 1347 873 1351
rect 405 1342 413 1346
rect -182 1331 -178 1339
rect -174 1331 -170 1339
rect 1106 1323 1114 1327
rect 1196 1323 1204 1327
rect 1372 1322 1380 1326
rect 1462 1322 1470 1326
rect 1106 1315 1114 1319
rect 1196 1315 1204 1319
rect 1372 1314 1380 1318
rect 1462 1314 1470 1318
rect 951 1310 959 1314
rect 865 1303 873 1307
rect 951 1302 959 1306
rect -113 1293 -105 1297
rect -23 1293 -15 1297
rect 153 1292 161 1296
rect 243 1292 251 1296
rect -113 1285 -105 1289
rect -23 1285 -15 1289
rect 153 1284 161 1288
rect 360 1289 368 1293
rect 865 1295 873 1299
rect 243 1284 251 1288
rect 360 1281 368 1285
rect 805 1283 813 1287
rect 397 1272 401 1280
rect 405 1272 409 1280
rect 805 1275 813 1279
rect 1106 1271 1114 1275
rect 1196 1271 1204 1275
rect 1372 1270 1380 1274
rect 1462 1270 1470 1274
rect 865 1260 873 1264
rect 951 1258 959 1262
rect 1106 1263 1114 1267
rect 1196 1263 1204 1267
rect 1372 1262 1380 1266
rect 1462 1262 1470 1266
rect 865 1252 873 1256
rect -172 1244 -164 1248
rect 951 1250 959 1254
rect -113 1241 -105 1245
rect -23 1241 -15 1245
rect 94 1243 102 1247
rect 153 1240 161 1244
rect -172 1236 -164 1240
rect 243 1240 251 1244
rect -113 1233 -105 1237
rect -23 1233 -15 1237
rect 94 1235 102 1239
rect 360 1237 368 1241
rect 153 1232 161 1236
rect 243 1232 251 1236
rect 360 1229 368 1233
rect 1041 1231 1045 1239
rect 1049 1231 1053 1239
rect 865 1208 873 1212
rect 865 1200 873 1204
rect -172 1192 -164 1196
rect 94 1191 102 1195
rect 1110 1193 1118 1197
rect 1200 1193 1208 1197
rect -172 1184 -164 1188
rect 94 1183 102 1187
rect 320 1183 324 1191
rect 328 1183 332 1191
rect 1376 1192 1384 1196
rect 1466 1192 1474 1196
rect 1110 1185 1118 1189
rect 1200 1185 1208 1189
rect 1376 1184 1384 1188
rect 1466 1184 1474 1188
rect 405 1162 413 1166
rect -117 1151 -109 1155
rect -27 1151 -19 1155
rect 149 1150 157 1154
rect 405 1154 413 1158
rect 239 1150 247 1154
rect -117 1143 -109 1147
rect -27 1143 -19 1147
rect 149 1142 157 1146
rect 239 1142 247 1146
rect 780 1143 784 1151
rect 788 1143 792 1151
rect 1051 1144 1059 1148
rect 1110 1141 1118 1145
rect 1200 1141 1208 1145
rect 1317 1143 1325 1147
rect 1376 1140 1384 1144
rect 1051 1136 1059 1140
rect 1466 1140 1474 1144
rect 491 1117 499 1121
rect 865 1122 873 1126
rect 1110 1133 1118 1137
rect 1200 1133 1208 1137
rect 1317 1135 1325 1139
rect 1376 1132 1384 1136
rect 1466 1132 1474 1136
rect 865 1114 873 1118
rect 405 1110 413 1114
rect 491 1109 499 1113
rect -117 1099 -109 1103
rect -27 1099 -19 1103
rect 149 1098 157 1102
rect 239 1098 247 1102
rect 405 1102 413 1106
rect -117 1091 -109 1095
rect -27 1091 -19 1095
rect 149 1090 157 1094
rect 239 1090 247 1094
rect 345 1090 353 1094
rect 345 1082 353 1086
rect 1051 1092 1059 1096
rect 1317 1091 1325 1095
rect 1051 1084 1059 1088
rect 951 1077 959 1081
rect 1317 1083 1325 1087
rect -182 1059 -178 1067
rect -174 1059 -170 1067
rect 405 1067 413 1071
rect 865 1070 873 1074
rect 951 1069 959 1073
rect 491 1065 499 1069
rect 405 1059 413 1063
rect 491 1057 499 1061
rect 865 1062 873 1066
rect 805 1050 813 1054
rect 1106 1051 1114 1055
rect 1196 1051 1204 1055
rect 1372 1050 1380 1054
rect 1462 1050 1470 1054
rect 805 1042 813 1046
rect 1106 1043 1114 1047
rect 1196 1043 1204 1047
rect 1372 1042 1380 1046
rect 1462 1042 1470 1046
rect -113 1021 -105 1025
rect -23 1021 -15 1025
rect 153 1020 161 1024
rect 243 1020 251 1024
rect 542 1023 546 1031
rect 550 1023 554 1031
rect 580 1023 584 1031
rect 588 1023 592 1031
rect 618 1023 622 1031
rect 626 1023 630 1031
rect 656 1023 660 1031
rect 664 1023 668 1031
rect 725 1024 729 1032
rect 733 1024 737 1032
rect 865 1027 873 1031
rect 951 1025 959 1029
rect -113 1013 -105 1017
rect -23 1013 -15 1017
rect 153 1012 161 1016
rect 243 1012 251 1016
rect 405 1015 413 1019
rect 405 1007 413 1011
rect 865 1019 873 1023
rect 951 1017 959 1021
rect 1106 999 1114 1003
rect 1196 999 1204 1003
rect 1372 998 1380 1002
rect 1462 998 1470 1002
rect 1106 991 1114 995
rect 1196 991 1204 995
rect 1372 990 1380 994
rect 1462 990 1470 994
rect -172 972 -164 976
rect -113 969 -105 973
rect -23 969 -15 973
rect 94 971 102 975
rect 865 975 873 979
rect 153 968 161 972
rect -172 964 -164 968
rect 243 968 251 972
rect -113 961 -105 965
rect -23 961 -15 965
rect 94 963 102 967
rect 725 967 729 975
rect 733 967 737 975
rect 153 960 161 964
rect 243 960 251 964
rect 360 954 368 958
rect 865 967 873 971
rect 1041 959 1045 967
rect 1049 959 1053 967
rect 360 946 368 950
rect 397 937 401 945
rect 405 937 409 945
rect -172 920 -164 924
rect 94 919 102 923
rect -172 912 -164 916
rect 94 911 102 915
rect 1110 921 1118 925
rect 1200 921 1208 925
rect 1376 920 1384 924
rect 1466 920 1474 924
rect 725 910 729 918
rect 733 910 737 918
rect 780 910 784 918
rect 788 910 792 918
rect 1110 913 1118 917
rect 1200 913 1208 917
rect 1376 912 1384 916
rect 1466 912 1474 916
rect 360 902 368 906
rect 360 894 368 898
rect -117 879 -109 883
rect -27 879 -19 883
rect 149 878 157 882
rect 865 889 873 893
rect 239 878 247 882
rect 865 881 873 885
rect -117 871 -109 875
rect -27 871 -19 875
rect 149 870 157 874
rect 239 870 247 874
rect 1051 872 1059 876
rect 1110 869 1118 873
rect 1200 869 1208 873
rect 1317 871 1325 875
rect 1376 868 1384 872
rect 1051 864 1059 868
rect 1466 868 1474 872
rect 320 848 324 856
rect 328 848 332 856
rect 725 853 729 861
rect 733 853 737 861
rect 1110 861 1118 865
rect 1200 861 1208 865
rect 1317 863 1325 867
rect 1376 860 1384 864
rect 1466 860 1474 864
rect 951 844 959 848
rect -117 827 -109 831
rect -27 827 -19 831
rect 149 826 157 830
rect 239 826 247 830
rect 865 837 873 841
rect 951 836 959 840
rect 405 827 413 831
rect -117 819 -109 823
rect 865 829 873 833
rect -27 819 -19 823
rect 149 818 157 822
rect 239 818 247 822
rect 405 819 413 823
rect 805 817 813 821
rect 1051 820 1059 824
rect 1317 819 1325 823
rect 805 809 813 813
rect 1051 812 1059 816
rect 1317 811 1325 815
rect -182 787 -178 795
rect -174 787 -170 795
rect 865 794 873 798
rect 951 792 959 796
rect 865 786 873 790
rect 491 782 499 786
rect 951 784 959 788
rect 405 775 413 779
rect 491 774 499 778
rect 1106 779 1114 783
rect 1196 779 1204 783
rect 1372 778 1380 782
rect 1462 778 1470 782
rect 405 767 413 771
rect 1106 771 1114 775
rect 1196 771 1204 775
rect 1372 770 1380 774
rect 1462 770 1470 774
rect -113 749 -105 753
rect -23 749 -15 753
rect 153 748 161 752
rect 345 755 353 759
rect 243 748 251 752
rect 345 747 353 751
rect -113 741 -105 745
rect -23 741 -15 745
rect 153 740 161 744
rect 243 740 251 744
rect 865 742 873 746
rect 405 732 413 736
rect 491 730 499 734
rect 865 734 873 738
rect 405 724 413 728
rect 1106 727 1114 731
rect 1196 727 1204 731
rect 1372 726 1380 730
rect 491 722 499 726
rect 1462 726 1470 730
rect 1106 719 1114 723
rect 1196 719 1204 723
rect 1372 718 1380 722
rect 1462 718 1470 722
rect -172 700 -164 704
rect -113 697 -105 701
rect -23 697 -15 701
rect 94 699 102 703
rect 153 696 161 700
rect -172 692 -164 696
rect 243 696 251 700
rect -113 689 -105 693
rect -23 689 -15 693
rect 94 691 102 695
rect 153 688 161 692
rect 243 688 251 692
rect 1041 687 1045 695
rect 1049 687 1053 695
rect 405 680 413 684
rect 780 677 784 685
rect 788 677 792 685
rect 405 672 413 676
rect 865 656 873 660
rect -172 648 -164 652
rect 94 647 102 651
rect 865 648 873 652
rect 1110 649 1118 653
rect 1200 649 1208 653
rect -172 640 -164 644
rect 1376 648 1384 652
rect 1466 648 1474 652
rect 94 639 102 643
rect 1110 641 1118 645
rect 1200 641 1208 645
rect 1376 640 1384 644
rect 1466 640 1474 644
rect 360 619 368 623
rect -117 607 -109 611
rect -27 607 -19 611
rect 149 606 157 610
rect 360 611 368 615
rect 951 611 959 615
rect 239 606 247 610
rect -117 599 -109 603
rect -27 599 -19 603
rect 149 598 157 602
rect 239 598 247 602
rect 397 602 401 610
rect 405 602 409 610
rect 865 604 873 608
rect 951 603 959 607
rect 865 596 873 600
rect 1051 600 1059 604
rect 1110 597 1118 601
rect 1200 597 1208 601
rect 1317 599 1325 603
rect 1376 596 1384 600
rect 1051 592 1059 596
rect 1466 596 1474 600
rect 805 584 813 588
rect 805 576 813 580
rect 1110 589 1118 593
rect 1200 589 1208 593
rect 1317 591 1325 595
rect 1376 588 1384 592
rect 1466 588 1474 592
rect 360 567 368 571
rect -117 555 -109 559
rect -27 555 -19 559
rect 149 554 157 558
rect 239 554 247 558
rect 360 559 368 563
rect 865 561 873 565
rect 951 559 959 563
rect 865 553 873 557
rect -117 547 -109 551
rect -27 547 -19 551
rect 149 546 157 550
rect 239 546 247 550
rect 951 551 959 555
rect 1051 548 1059 552
rect 1317 547 1325 551
rect 1051 540 1059 544
rect 1317 539 1325 543
rect -182 515 -178 523
rect -174 515 -170 523
rect 320 513 324 521
rect 328 513 332 521
rect 865 509 873 513
rect 1106 507 1114 511
rect 1196 507 1204 511
rect 865 501 873 505
rect 1372 506 1380 510
rect 1462 506 1470 510
rect 1106 499 1114 503
rect 1196 499 1204 503
rect 1372 498 1380 502
rect 1462 498 1470 502
rect 405 492 413 496
rect 405 484 413 488
rect -113 477 -105 481
rect -23 477 -15 481
rect 153 476 161 480
rect 243 476 251 480
rect -113 469 -105 473
rect -23 469 -15 473
rect 153 468 161 472
rect 243 468 251 472
rect 1106 455 1114 459
rect 1196 455 1204 459
rect 1372 454 1380 458
rect 1462 454 1470 458
rect 491 447 499 451
rect 1106 447 1114 451
rect 1196 447 1204 451
rect 405 440 413 444
rect 1372 446 1380 450
rect 1462 446 1470 450
rect 491 439 499 443
rect -172 428 -164 432
rect -113 425 -105 429
rect -23 425 -15 429
rect 94 427 102 431
rect 153 424 161 428
rect -172 420 -164 424
rect 243 424 251 428
rect 405 432 413 436
rect -113 417 -105 421
rect -23 417 -15 421
rect 94 419 102 423
rect 153 416 161 420
rect 243 416 251 420
rect 345 420 353 424
rect 345 412 353 416
rect 1041 415 1045 423
rect 1049 415 1053 423
rect 405 397 413 401
rect 491 395 499 399
rect 405 389 413 393
rect 491 387 499 391
rect -172 376 -164 380
rect 94 375 102 379
rect 1110 377 1118 381
rect 1200 377 1208 381
rect -172 368 -164 372
rect 1376 376 1384 380
rect 1466 376 1474 380
rect 94 367 102 371
rect 1110 369 1118 373
rect 1200 369 1208 373
rect 1376 368 1384 372
rect 1466 368 1474 372
rect 405 345 413 349
rect -117 335 -109 339
rect -27 335 -19 339
rect 149 334 157 338
rect 239 334 247 338
rect 405 337 413 341
rect -117 327 -109 331
rect -27 327 -19 331
rect 149 326 157 330
rect 239 326 247 330
rect 1051 328 1059 332
rect 1110 325 1118 329
rect 1200 325 1208 329
rect 1317 327 1325 331
rect 1376 324 1384 328
rect 1051 320 1059 324
rect 1466 324 1474 328
rect 1110 317 1118 321
rect 1200 317 1208 321
rect 1317 319 1325 323
rect 1376 316 1384 320
rect 1466 316 1474 320
rect -117 283 -109 287
rect -27 283 -19 287
rect 149 282 157 286
rect 239 282 247 286
rect 360 284 368 288
rect -117 275 -109 279
rect -27 275 -19 279
rect 149 274 157 278
rect 239 274 247 278
rect 360 276 368 280
rect 1051 276 1059 280
rect 1317 275 1325 279
rect 397 267 401 275
rect 405 267 409 275
rect 1051 268 1059 272
rect 1317 267 1325 271
rect -182 243 -178 251
rect -174 243 -170 251
rect 360 232 368 236
rect 360 224 368 228
rect -113 205 -105 209
rect -23 205 -15 209
rect 153 204 161 208
rect 243 204 251 208
rect -113 197 -105 201
rect -23 197 -15 201
rect 153 196 161 200
rect 243 196 251 200
rect -172 156 -164 160
rect -113 153 -105 157
rect -23 153 -15 157
rect 94 155 102 159
rect 153 152 161 156
rect -172 148 -164 152
rect 243 152 251 156
rect -113 145 -105 149
rect -23 145 -15 149
rect 94 147 102 151
rect 153 144 161 148
rect 243 144 251 148
rect -172 104 -164 108
rect 94 103 102 107
rect -172 96 -164 100
rect 94 95 102 99
rect -117 63 -109 67
rect -27 63 -19 67
rect 149 62 157 66
rect 239 62 247 66
rect -117 55 -109 59
rect -27 55 -19 59
rect 149 54 157 58
rect 239 54 247 58
rect -117 11 -109 15
rect -27 11 -19 15
rect 149 10 157 14
rect 239 10 247 14
rect -117 3 -109 7
rect -27 3 -19 7
rect 149 2 157 6
rect 239 2 247 6
rect -182 -29 -178 -21
rect -174 -29 -170 -21
rect -113 -67 -105 -63
rect -23 -67 -15 -63
rect 153 -68 161 -64
rect 243 -68 251 -64
rect -113 -75 -105 -71
rect -23 -75 -15 -71
rect 153 -76 161 -72
rect 243 -76 251 -72
rect -172 -116 -164 -112
rect -113 -119 -105 -115
rect -23 -119 -15 -115
rect 94 -117 102 -113
rect 153 -120 161 -116
rect -172 -124 -164 -120
rect 243 -120 251 -116
rect -113 -127 -105 -123
rect -23 -127 -15 -123
rect 94 -125 102 -121
rect 153 -128 161 -124
rect 243 -128 251 -124
rect -172 -168 -164 -164
rect 94 -169 102 -165
rect -172 -176 -164 -172
rect 94 -177 102 -173
<< polysilicon >>
rect -127 1966 -125 1970
rect -37 1966 -35 1970
rect -130 1964 -117 1966
rect -109 1964 -106 1966
rect -40 1964 -27 1966
rect -19 1964 -16 1966
rect 139 1965 141 1969
rect 229 1965 231 1969
rect 136 1963 149 1965
rect 157 1963 160 1965
rect 226 1963 239 1965
rect 247 1963 250 1965
rect -150 1948 -148 1954
rect -60 1948 -58 1954
rect -166 1946 -163 1948
rect -155 1946 -145 1948
rect -76 1946 -73 1948
rect -65 1946 -55 1948
rect 116 1947 118 1953
rect 206 1947 208 1953
rect 100 1945 103 1947
rect 111 1945 121 1947
rect 190 1945 193 1947
rect 201 1945 211 1947
rect -151 1938 -141 1940
rect -133 1938 -130 1940
rect -61 1938 -51 1940
rect -43 1938 -40 1940
rect -147 1929 -145 1938
rect -57 1929 -55 1938
rect 115 1937 125 1939
rect 133 1937 136 1939
rect 205 1937 215 1939
rect 223 1937 226 1939
rect 119 1928 121 1937
rect 209 1928 211 1937
rect -130 1912 -117 1914
rect -109 1912 -106 1914
rect -40 1912 -27 1914
rect -19 1912 -16 1914
rect -127 1908 -125 1912
rect -37 1908 -35 1912
rect 136 1911 149 1913
rect 157 1911 160 1913
rect 226 1911 239 1913
rect 247 1911 250 1913
rect 139 1907 141 1911
rect 229 1907 231 1911
rect -177 1883 -175 1886
rect -177 1867 -175 1875
rect -185 1865 -175 1867
rect -177 1863 -175 1865
rect -177 1852 -175 1855
rect -123 1836 -121 1840
rect -33 1836 -31 1840
rect -126 1834 -113 1836
rect -105 1834 -102 1836
rect -36 1834 -23 1836
rect -15 1834 -12 1836
rect 143 1835 145 1839
rect 233 1835 235 1839
rect 140 1833 153 1835
rect 161 1833 164 1835
rect 230 1833 243 1835
rect 251 1833 254 1835
rect -146 1818 -144 1824
rect -56 1818 -54 1824
rect -162 1816 -159 1818
rect -151 1816 -141 1818
rect -72 1816 -69 1818
rect -61 1816 -51 1818
rect 120 1817 122 1823
rect 210 1817 212 1823
rect 104 1815 107 1817
rect 115 1815 125 1817
rect 194 1815 197 1817
rect 205 1815 215 1817
rect -147 1808 -137 1810
rect -129 1808 -126 1810
rect -57 1808 -47 1810
rect -39 1808 -36 1810
rect -143 1799 -141 1808
rect -53 1799 -51 1808
rect 119 1807 129 1809
rect 137 1807 140 1809
rect 209 1807 219 1809
rect 227 1807 230 1809
rect 123 1798 125 1807
rect 213 1798 215 1807
rect -182 1787 -180 1791
rect -185 1785 -172 1787
rect -164 1785 -161 1787
rect 84 1786 86 1790
rect 81 1784 94 1786
rect 102 1784 105 1786
rect -126 1782 -113 1784
rect -105 1782 -102 1784
rect -36 1782 -23 1784
rect -15 1782 -12 1784
rect -123 1778 -121 1782
rect -205 1769 -203 1775
rect -33 1778 -31 1782
rect 140 1781 153 1783
rect 161 1781 164 1783
rect 230 1781 243 1783
rect 251 1781 254 1783
rect 143 1777 145 1781
rect -221 1767 -218 1769
rect -210 1767 -200 1769
rect 61 1768 63 1774
rect 233 1777 235 1781
rect 45 1766 48 1768
rect 56 1766 66 1768
rect -206 1759 -196 1761
rect -188 1759 -185 1761
rect -202 1750 -200 1759
rect 60 1758 70 1760
rect 78 1758 81 1760
rect 64 1749 66 1758
rect -185 1733 -172 1735
rect -164 1733 -161 1735
rect -182 1729 -180 1733
rect 81 1732 94 1734
rect 102 1732 105 1734
rect 84 1728 86 1732
rect -127 1694 -125 1698
rect -37 1694 -35 1698
rect -130 1692 -117 1694
rect -109 1692 -106 1694
rect -40 1692 -27 1694
rect -19 1692 -16 1694
rect 139 1693 141 1697
rect 229 1693 231 1697
rect 136 1691 149 1693
rect 157 1691 160 1693
rect 226 1691 239 1693
rect 247 1691 250 1693
rect -150 1676 -148 1682
rect -60 1676 -58 1682
rect -166 1674 -163 1676
rect -155 1674 -145 1676
rect -76 1674 -73 1676
rect -65 1674 -55 1676
rect 116 1675 118 1681
rect 206 1675 208 1681
rect 100 1673 103 1675
rect 111 1673 121 1675
rect 190 1673 193 1675
rect 201 1673 211 1675
rect -151 1666 -141 1668
rect -133 1666 -130 1668
rect -61 1666 -51 1668
rect -43 1666 -40 1668
rect -147 1657 -145 1666
rect -57 1657 -55 1666
rect 115 1665 125 1667
rect 133 1665 136 1667
rect 205 1665 215 1667
rect 223 1665 226 1667
rect 119 1656 121 1665
rect 209 1656 211 1665
rect -130 1640 -117 1642
rect -109 1640 -106 1642
rect -40 1640 -27 1642
rect -19 1640 -16 1642
rect -127 1636 -125 1640
rect -37 1636 -35 1640
rect 136 1639 149 1641
rect 157 1639 160 1641
rect 226 1639 239 1641
rect 247 1639 250 1641
rect 139 1635 141 1639
rect 229 1635 231 1639
rect -177 1611 -175 1614
rect -177 1595 -175 1603
rect -185 1593 -175 1595
rect 1096 1594 1098 1598
rect 1186 1594 1188 1598
rect -177 1591 -175 1593
rect 1093 1592 1106 1594
rect 1114 1592 1117 1594
rect 1183 1592 1196 1594
rect 1204 1592 1207 1594
rect 1362 1593 1364 1597
rect 1452 1593 1454 1597
rect 1359 1591 1372 1593
rect 1380 1591 1383 1593
rect 1449 1591 1462 1593
rect 1470 1591 1473 1593
rect -177 1580 -175 1583
rect 1073 1576 1075 1582
rect 1163 1576 1165 1582
rect 1057 1574 1060 1576
rect 1068 1574 1078 1576
rect 1147 1574 1150 1576
rect 1158 1574 1168 1576
rect 1339 1575 1341 1581
rect 1429 1575 1431 1581
rect 1323 1573 1326 1575
rect 1334 1573 1344 1575
rect 1413 1573 1416 1575
rect 1424 1573 1434 1575
rect -123 1564 -121 1568
rect -33 1564 -31 1568
rect -126 1562 -113 1564
rect -105 1562 -102 1564
rect -36 1562 -23 1564
rect -15 1562 -12 1564
rect 143 1563 145 1567
rect 233 1563 235 1567
rect 1072 1566 1082 1568
rect 1090 1566 1093 1568
rect 1162 1566 1172 1568
rect 1180 1566 1183 1568
rect 140 1561 153 1563
rect 161 1561 164 1563
rect 230 1561 243 1563
rect 251 1561 254 1563
rect 1076 1557 1078 1566
rect 1166 1557 1168 1566
rect 1338 1565 1348 1567
rect 1356 1565 1359 1567
rect 1428 1565 1438 1567
rect 1446 1565 1449 1567
rect -146 1546 -144 1552
rect -56 1546 -54 1552
rect 1342 1556 1344 1565
rect 1432 1556 1434 1565
rect -162 1544 -159 1546
rect -151 1544 -141 1546
rect -72 1544 -69 1546
rect -61 1544 -51 1546
rect 120 1545 122 1551
rect 210 1545 212 1551
rect 104 1543 107 1545
rect 115 1543 125 1545
rect 194 1543 197 1545
rect 205 1543 215 1545
rect 1093 1540 1106 1542
rect 1114 1540 1117 1542
rect 1183 1540 1196 1542
rect 1204 1540 1207 1542
rect -147 1536 -137 1538
rect -129 1536 -126 1538
rect -57 1536 -47 1538
rect -39 1536 -36 1538
rect -143 1527 -141 1536
rect -53 1527 -51 1536
rect 119 1535 129 1537
rect 137 1535 140 1537
rect 209 1535 219 1537
rect 227 1535 230 1537
rect 1096 1536 1098 1540
rect 123 1526 125 1535
rect 213 1526 215 1535
rect 1186 1536 1188 1540
rect 1359 1539 1372 1541
rect 1380 1539 1383 1541
rect 1449 1539 1462 1541
rect 1470 1539 1473 1541
rect 1362 1535 1364 1539
rect 1452 1535 1454 1539
rect 325 1526 327 1529
rect -182 1515 -180 1519
rect -185 1513 -172 1515
rect -164 1513 -161 1515
rect 84 1514 86 1518
rect 81 1512 94 1514
rect 102 1512 105 1514
rect -126 1510 -113 1512
rect -105 1510 -102 1512
rect -36 1510 -23 1512
rect -15 1510 -12 1512
rect -123 1506 -121 1510
rect -205 1497 -203 1503
rect -33 1506 -31 1510
rect 140 1509 153 1511
rect 161 1509 164 1511
rect 230 1509 243 1511
rect 251 1509 254 1511
rect 143 1505 145 1509
rect -221 1495 -218 1497
rect -210 1495 -200 1497
rect 61 1496 63 1502
rect 233 1505 235 1509
rect 325 1510 327 1518
rect 1046 1511 1048 1514
rect 317 1508 327 1510
rect 325 1506 327 1508
rect 45 1494 48 1496
rect 56 1494 66 1496
rect 325 1495 327 1498
rect 395 1496 397 1500
rect 392 1494 405 1496
rect 413 1494 416 1496
rect 1046 1495 1048 1503
rect 1038 1493 1048 1495
rect 1046 1491 1048 1493
rect -206 1487 -196 1489
rect -188 1487 -185 1489
rect -202 1478 -200 1487
rect 60 1486 70 1488
rect 78 1486 81 1488
rect 64 1477 66 1486
rect 372 1478 374 1484
rect 1046 1480 1048 1483
rect 356 1476 359 1478
rect 367 1476 377 1478
rect 371 1468 381 1470
rect 389 1468 392 1470
rect -185 1461 -172 1463
rect -164 1461 -161 1463
rect -182 1457 -180 1461
rect 81 1460 94 1462
rect 102 1460 105 1462
rect 84 1456 86 1460
rect 375 1459 377 1468
rect 1100 1464 1102 1468
rect 1190 1464 1192 1468
rect 1097 1462 1110 1464
rect 1118 1462 1121 1464
rect 1187 1462 1200 1464
rect 1208 1462 1211 1464
rect 1366 1463 1368 1467
rect 1456 1463 1458 1467
rect 1363 1461 1376 1463
rect 1384 1461 1387 1463
rect 1453 1461 1466 1463
rect 1474 1461 1477 1463
rect 481 1451 483 1455
rect 478 1449 491 1451
rect 499 1449 502 1451
rect 1077 1446 1079 1452
rect 1167 1446 1169 1452
rect 1061 1444 1064 1446
rect 1072 1444 1082 1446
rect 1151 1444 1154 1446
rect 1162 1444 1172 1446
rect 1343 1445 1345 1451
rect 1433 1445 1435 1451
rect 392 1442 405 1444
rect 413 1442 416 1444
rect 1327 1443 1330 1445
rect 1338 1443 1348 1445
rect 1417 1443 1420 1445
rect 1428 1443 1438 1445
rect 395 1438 397 1442
rect 458 1433 460 1439
rect 1076 1436 1086 1438
rect 1094 1436 1097 1438
rect 1166 1436 1176 1438
rect 1184 1436 1187 1438
rect -127 1422 -125 1426
rect -37 1422 -35 1426
rect -130 1420 -117 1422
rect -109 1420 -106 1422
rect -40 1420 -27 1422
rect -19 1420 -16 1422
rect 139 1421 141 1425
rect 229 1421 231 1425
rect 335 1424 337 1432
rect 442 1431 445 1433
rect 453 1431 463 1433
rect 1080 1427 1082 1436
rect 1170 1427 1172 1436
rect 1342 1435 1352 1437
rect 1360 1435 1363 1437
rect 1432 1435 1442 1437
rect 1450 1435 1453 1437
rect 322 1422 325 1424
rect 333 1422 345 1424
rect 353 1422 356 1424
rect 457 1423 467 1425
rect 475 1423 478 1425
rect 1346 1426 1348 1435
rect 1436 1426 1438 1435
rect 136 1419 149 1421
rect 157 1419 160 1421
rect 226 1419 239 1421
rect 247 1419 250 1421
rect 461 1414 463 1423
rect 1041 1415 1043 1419
rect -150 1404 -148 1410
rect -60 1404 -58 1410
rect 1038 1413 1051 1415
rect 1059 1413 1062 1415
rect 1307 1414 1309 1418
rect 1304 1412 1317 1414
rect 1325 1412 1328 1414
rect -166 1402 -163 1404
rect -155 1402 -145 1404
rect -76 1402 -73 1404
rect -65 1402 -55 1404
rect 116 1403 118 1409
rect 206 1403 208 1409
rect 1097 1410 1110 1412
rect 1118 1410 1121 1412
rect 1187 1410 1200 1412
rect 1208 1410 1211 1412
rect 100 1401 103 1403
rect 111 1401 121 1403
rect 190 1401 193 1403
rect 201 1401 211 1403
rect 395 1401 397 1405
rect 392 1399 405 1401
rect 413 1399 416 1401
rect 1100 1406 1102 1410
rect -151 1394 -141 1396
rect -133 1394 -130 1396
rect -61 1394 -51 1396
rect -43 1394 -40 1396
rect -147 1385 -145 1394
rect -57 1385 -55 1394
rect 115 1393 125 1395
rect 133 1393 136 1395
rect 205 1393 215 1395
rect 223 1393 226 1395
rect 478 1397 491 1399
rect 499 1397 502 1399
rect 1018 1397 1020 1403
rect 1190 1406 1192 1410
rect 1363 1409 1376 1411
rect 1384 1409 1387 1411
rect 1453 1409 1466 1411
rect 1474 1409 1477 1411
rect 1366 1405 1368 1409
rect 481 1393 483 1397
rect 119 1384 121 1393
rect 209 1384 211 1393
rect 1002 1395 1005 1397
rect 1013 1395 1023 1397
rect 1284 1396 1286 1402
rect 1456 1405 1458 1409
rect 1268 1394 1271 1396
rect 1279 1394 1289 1396
rect 372 1383 374 1389
rect 1017 1387 1027 1389
rect 1035 1387 1038 1389
rect 785 1384 787 1387
rect 356 1381 359 1383
rect 367 1381 377 1383
rect 1021 1378 1023 1387
rect 1283 1386 1293 1388
rect 1301 1386 1304 1388
rect -130 1368 -117 1370
rect -109 1368 -106 1370
rect -40 1368 -27 1370
rect -19 1368 -16 1370
rect 371 1373 381 1375
rect 389 1373 392 1375
rect -127 1364 -125 1368
rect -37 1364 -35 1368
rect 136 1367 149 1369
rect 157 1367 160 1369
rect 226 1367 239 1369
rect 247 1367 250 1369
rect 139 1363 141 1367
rect 229 1363 231 1367
rect 375 1364 377 1373
rect 785 1368 787 1376
rect 1287 1377 1289 1386
rect 777 1366 787 1368
rect 785 1364 787 1366
rect 1038 1361 1051 1363
rect 1059 1361 1062 1363
rect 785 1353 787 1356
rect 855 1354 857 1358
rect 1041 1357 1043 1361
rect 1304 1360 1317 1362
rect 1325 1360 1328 1362
rect 852 1352 865 1354
rect 873 1352 876 1354
rect 1307 1356 1309 1360
rect 392 1347 405 1349
rect 413 1347 416 1349
rect 395 1343 397 1347
rect -177 1339 -175 1342
rect 832 1336 834 1342
rect 816 1334 819 1336
rect 827 1334 837 1336
rect -177 1323 -175 1331
rect 831 1326 841 1328
rect 849 1326 852 1328
rect -185 1321 -175 1323
rect -177 1319 -175 1321
rect 835 1317 837 1326
rect 1096 1322 1098 1326
rect 1186 1322 1188 1326
rect 1093 1320 1106 1322
rect 1114 1320 1117 1322
rect 1183 1320 1196 1322
rect 1204 1320 1207 1322
rect 1362 1321 1364 1325
rect 1452 1321 1454 1325
rect 1359 1319 1372 1321
rect 1380 1319 1383 1321
rect 1449 1319 1462 1321
rect 1470 1319 1473 1321
rect -177 1308 -175 1311
rect 941 1309 943 1313
rect 938 1307 951 1309
rect 959 1307 962 1309
rect 1073 1304 1075 1310
rect 1163 1304 1165 1310
rect 1057 1302 1060 1304
rect 1068 1302 1078 1304
rect 1147 1302 1150 1304
rect 1158 1302 1168 1304
rect 1339 1303 1341 1309
rect 1429 1303 1431 1309
rect 852 1300 865 1302
rect 873 1300 876 1302
rect 1323 1301 1326 1303
rect 1334 1301 1344 1303
rect 1413 1301 1416 1303
rect 1424 1301 1434 1303
rect -123 1292 -121 1296
rect -33 1292 -31 1296
rect -126 1290 -113 1292
rect -105 1290 -102 1292
rect -36 1290 -23 1292
rect -15 1290 -12 1292
rect 143 1291 145 1295
rect 855 1296 857 1300
rect 233 1291 235 1295
rect 140 1289 153 1291
rect 161 1289 164 1291
rect 230 1289 243 1291
rect 251 1289 254 1291
rect 350 1288 352 1292
rect 918 1291 920 1297
rect 1072 1294 1082 1296
rect 1090 1294 1093 1296
rect 1162 1294 1172 1296
rect 1180 1294 1183 1296
rect 347 1286 360 1288
rect 368 1286 371 1288
rect -146 1274 -144 1280
rect -56 1274 -54 1280
rect 402 1280 404 1283
rect 795 1282 797 1290
rect 902 1289 905 1291
rect 913 1289 923 1291
rect 1076 1285 1078 1294
rect 1166 1285 1168 1294
rect 1338 1293 1348 1295
rect 1356 1293 1359 1295
rect 1428 1293 1438 1295
rect 1446 1293 1449 1295
rect 782 1280 785 1282
rect 793 1280 805 1282
rect 813 1280 816 1282
rect 917 1281 927 1283
rect 935 1281 938 1283
rect 1342 1284 1344 1293
rect 1432 1284 1434 1293
rect -162 1272 -159 1274
rect -151 1272 -141 1274
rect -72 1272 -69 1274
rect -61 1272 -51 1274
rect 120 1273 122 1279
rect 210 1273 212 1279
rect 104 1271 107 1273
rect 115 1271 125 1273
rect 194 1271 197 1273
rect 205 1271 215 1273
rect 327 1270 329 1276
rect 921 1272 923 1281
rect 311 1268 314 1270
rect 322 1268 332 1270
rect -147 1264 -137 1266
rect -129 1264 -126 1266
rect -57 1264 -47 1266
rect -39 1264 -36 1266
rect -143 1255 -141 1264
rect -53 1255 -51 1264
rect 119 1263 129 1265
rect 137 1263 140 1265
rect 209 1263 219 1265
rect 227 1263 230 1265
rect 123 1254 125 1263
rect 213 1254 215 1263
rect 326 1260 336 1262
rect 344 1260 347 1262
rect 402 1264 404 1272
rect 1093 1268 1106 1270
rect 1114 1268 1117 1270
rect 1183 1268 1196 1270
rect 1204 1268 1207 1270
rect 394 1262 404 1264
rect 1096 1264 1098 1268
rect 402 1260 404 1262
rect 330 1251 332 1260
rect 855 1259 857 1263
rect 852 1257 865 1259
rect 873 1257 876 1259
rect 1186 1264 1188 1268
rect 1359 1267 1372 1269
rect 1380 1267 1383 1269
rect 1449 1267 1462 1269
rect 1470 1267 1473 1269
rect 1362 1263 1364 1267
rect 1452 1263 1454 1267
rect 938 1255 951 1257
rect 959 1255 962 1257
rect -182 1243 -180 1247
rect 402 1249 404 1252
rect 941 1251 943 1255
rect -185 1241 -172 1243
rect -164 1241 -161 1243
rect 84 1242 86 1246
rect 81 1240 94 1242
rect 102 1240 105 1242
rect -126 1238 -113 1240
rect -105 1238 -102 1240
rect -36 1238 -23 1240
rect -15 1238 -12 1240
rect 832 1241 834 1247
rect -123 1234 -121 1238
rect -205 1225 -203 1231
rect -33 1234 -31 1238
rect 140 1237 153 1239
rect 161 1237 164 1239
rect 230 1237 243 1239
rect 251 1237 254 1239
rect 816 1239 819 1241
rect 827 1239 837 1241
rect 1046 1239 1048 1242
rect 143 1233 145 1237
rect -221 1223 -218 1225
rect -210 1223 -200 1225
rect 61 1224 63 1230
rect 233 1233 235 1237
rect 347 1234 360 1236
rect 368 1234 371 1236
rect 350 1230 352 1234
rect 831 1231 841 1233
rect 849 1231 852 1233
rect 45 1222 48 1224
rect 56 1222 66 1224
rect 835 1222 837 1231
rect 1046 1223 1048 1231
rect 1038 1221 1048 1223
rect 1046 1219 1048 1221
rect -206 1215 -196 1217
rect -188 1215 -185 1217
rect -202 1206 -200 1215
rect 60 1214 70 1216
rect 78 1214 81 1216
rect 64 1205 66 1214
rect 1046 1208 1048 1211
rect 852 1205 865 1207
rect 873 1205 876 1207
rect 855 1201 857 1205
rect 325 1191 327 1194
rect 1100 1192 1102 1196
rect 1190 1192 1192 1196
rect -185 1189 -172 1191
rect -164 1189 -161 1191
rect -182 1185 -180 1189
rect 81 1188 94 1190
rect 102 1188 105 1190
rect 84 1184 86 1188
rect 1097 1190 1110 1192
rect 1118 1190 1121 1192
rect 1187 1190 1200 1192
rect 1208 1190 1211 1192
rect 1366 1191 1368 1195
rect 1456 1191 1458 1195
rect 1363 1189 1376 1191
rect 1384 1189 1387 1191
rect 1453 1189 1466 1191
rect 1474 1189 1477 1191
rect 325 1175 327 1183
rect 317 1173 327 1175
rect 1077 1174 1079 1180
rect 1167 1174 1169 1180
rect 325 1171 327 1173
rect 1061 1172 1064 1174
rect 1072 1172 1082 1174
rect 1151 1172 1154 1174
rect 1162 1172 1172 1174
rect 1343 1173 1345 1179
rect 1433 1173 1435 1179
rect 1327 1171 1330 1173
rect 1338 1171 1348 1173
rect 1417 1171 1420 1173
rect 1428 1171 1438 1173
rect 325 1160 327 1163
rect 395 1161 397 1165
rect 1076 1164 1086 1166
rect 1094 1164 1097 1166
rect 1166 1164 1176 1166
rect 1184 1164 1187 1166
rect 392 1159 405 1161
rect 413 1159 416 1161
rect -127 1150 -125 1154
rect -37 1150 -35 1154
rect -130 1148 -117 1150
rect -109 1148 -106 1150
rect -40 1148 -27 1150
rect -19 1148 -16 1150
rect 139 1149 141 1153
rect 1080 1155 1082 1164
rect 1170 1155 1172 1164
rect 1342 1163 1352 1165
rect 1360 1163 1363 1165
rect 1432 1163 1442 1165
rect 1450 1163 1453 1165
rect 229 1149 231 1153
rect 785 1151 787 1154
rect 1346 1154 1348 1163
rect 1436 1154 1438 1163
rect 136 1147 149 1149
rect 157 1147 160 1149
rect 226 1147 239 1149
rect 247 1147 250 1149
rect 372 1143 374 1149
rect 1041 1143 1043 1147
rect 356 1141 359 1143
rect 367 1141 377 1143
rect -150 1132 -148 1138
rect -60 1132 -58 1138
rect -166 1130 -163 1132
rect -155 1130 -145 1132
rect -76 1130 -73 1132
rect -65 1130 -55 1132
rect 116 1131 118 1137
rect 206 1131 208 1137
rect 371 1133 381 1135
rect 389 1133 392 1135
rect 100 1129 103 1131
rect 111 1129 121 1131
rect 190 1129 193 1131
rect 201 1129 211 1131
rect 375 1124 377 1133
rect 785 1135 787 1143
rect 1038 1141 1051 1143
rect 1059 1141 1062 1143
rect 1307 1142 1309 1146
rect 1304 1140 1317 1142
rect 1325 1140 1328 1142
rect 1097 1138 1110 1140
rect 1118 1138 1121 1140
rect 1187 1138 1200 1140
rect 1208 1138 1211 1140
rect 777 1133 787 1135
rect 785 1131 787 1133
rect 1100 1134 1102 1138
rect -151 1122 -141 1124
rect -133 1122 -130 1124
rect -61 1122 -51 1124
rect -43 1122 -40 1124
rect -147 1113 -145 1122
rect -57 1113 -55 1122
rect 115 1121 125 1123
rect 133 1121 136 1123
rect 205 1121 215 1123
rect 223 1121 226 1123
rect 119 1112 121 1121
rect 209 1112 211 1121
rect 481 1116 483 1120
rect 785 1120 787 1123
rect 855 1121 857 1125
rect 1018 1125 1020 1131
rect 1190 1134 1192 1138
rect 1363 1137 1376 1139
rect 1384 1137 1387 1139
rect 1453 1137 1466 1139
rect 1474 1137 1477 1139
rect 1366 1133 1368 1137
rect 1002 1123 1005 1125
rect 1013 1123 1023 1125
rect 1284 1124 1286 1130
rect 1456 1133 1458 1137
rect 1268 1122 1271 1124
rect 1279 1122 1289 1124
rect 852 1119 865 1121
rect 873 1119 876 1121
rect 478 1114 491 1116
rect 499 1114 502 1116
rect 1017 1115 1027 1117
rect 1035 1115 1038 1117
rect 392 1107 405 1109
rect 413 1107 416 1109
rect 395 1103 397 1107
rect -130 1096 -117 1098
rect -109 1096 -106 1098
rect -40 1096 -27 1098
rect -19 1096 -16 1098
rect 458 1098 460 1104
rect 832 1103 834 1109
rect 1021 1106 1023 1115
rect 1283 1114 1293 1116
rect 1301 1114 1304 1116
rect 816 1101 819 1103
rect 827 1101 837 1103
rect 1287 1105 1289 1114
rect -127 1092 -125 1096
rect -37 1092 -35 1096
rect 136 1095 149 1097
rect 157 1095 160 1097
rect 226 1095 239 1097
rect 247 1095 250 1097
rect 139 1091 141 1095
rect 229 1091 231 1095
rect 335 1089 337 1097
rect 442 1096 445 1098
rect 453 1096 463 1098
rect 831 1093 841 1095
rect 849 1093 852 1095
rect 322 1087 325 1089
rect 333 1087 345 1089
rect 353 1087 356 1089
rect 457 1088 467 1090
rect 475 1088 478 1090
rect 461 1079 463 1088
rect 835 1084 837 1093
rect 1038 1089 1051 1091
rect 1059 1089 1062 1091
rect 1041 1085 1043 1089
rect 1304 1088 1317 1090
rect 1325 1088 1328 1090
rect 1307 1084 1309 1088
rect 941 1076 943 1080
rect 938 1074 951 1076
rect 959 1074 962 1076
rect -177 1067 -175 1070
rect 395 1066 397 1070
rect 392 1064 405 1066
rect 413 1064 416 1066
rect 852 1067 865 1069
rect 873 1067 876 1069
rect 478 1062 491 1064
rect 499 1062 502 1064
rect 855 1063 857 1067
rect -177 1051 -175 1059
rect 481 1058 483 1062
rect 918 1058 920 1064
rect -185 1049 -175 1051
rect -177 1047 -175 1049
rect 372 1048 374 1054
rect 795 1049 797 1057
rect 902 1056 905 1058
rect 913 1056 923 1058
rect 1096 1050 1098 1054
rect 1186 1050 1188 1054
rect 356 1046 359 1048
rect 367 1046 377 1048
rect 782 1047 785 1049
rect 793 1047 805 1049
rect 813 1047 816 1049
rect 917 1048 927 1050
rect 935 1048 938 1050
rect 1093 1048 1106 1050
rect 1114 1048 1117 1050
rect 1183 1048 1196 1050
rect 1204 1048 1207 1050
rect 1362 1049 1364 1053
rect 1452 1049 1454 1053
rect -177 1036 -175 1039
rect 371 1038 381 1040
rect 389 1038 392 1040
rect 921 1039 923 1048
rect 1359 1047 1372 1049
rect 1380 1047 1383 1049
rect 1449 1047 1462 1049
rect 1470 1047 1473 1049
rect 375 1029 377 1038
rect 547 1031 549 1034
rect 585 1031 587 1034
rect 623 1031 625 1034
rect 661 1031 663 1034
rect 730 1032 732 1035
rect -123 1020 -121 1024
rect -33 1020 -31 1024
rect -126 1018 -113 1020
rect -105 1018 -102 1020
rect -36 1018 -23 1020
rect -15 1018 -12 1020
rect 143 1019 145 1023
rect 233 1019 235 1023
rect 1073 1032 1075 1038
rect 1163 1032 1165 1038
rect 855 1026 857 1030
rect 1057 1030 1060 1032
rect 1068 1030 1078 1032
rect 1147 1030 1150 1032
rect 1158 1030 1168 1032
rect 1339 1031 1341 1037
rect 1429 1031 1431 1037
rect 1323 1029 1326 1031
rect 1334 1029 1344 1031
rect 1413 1029 1416 1031
rect 1424 1029 1434 1031
rect 852 1024 865 1026
rect 873 1024 876 1026
rect 140 1017 153 1019
rect 161 1017 164 1019
rect 230 1017 243 1019
rect 251 1017 254 1019
rect 392 1012 405 1014
rect 413 1012 416 1014
rect 547 1015 549 1023
rect 543 1013 549 1015
rect -146 1002 -144 1008
rect -56 1002 -54 1008
rect 395 1008 397 1012
rect -162 1000 -159 1002
rect -151 1000 -141 1002
rect -72 1000 -69 1002
rect -61 1000 -51 1002
rect 120 1001 122 1007
rect 210 1001 212 1007
rect 547 1010 549 1013
rect 585 1015 587 1023
rect 581 1013 587 1015
rect 585 1010 587 1013
rect 623 1015 625 1023
rect 619 1013 625 1015
rect 623 1010 625 1013
rect 661 1015 663 1023
rect 657 1013 663 1015
rect 730 1016 732 1024
rect 938 1022 951 1024
rect 959 1022 962 1024
rect 1072 1022 1082 1024
rect 1090 1022 1093 1024
rect 1162 1022 1172 1024
rect 1180 1022 1183 1024
rect 941 1018 943 1022
rect 722 1014 732 1016
rect 661 1010 663 1013
rect 730 1012 732 1014
rect 832 1008 834 1014
rect 1076 1013 1078 1022
rect 1166 1013 1168 1022
rect 1338 1021 1348 1023
rect 1356 1021 1359 1023
rect 1428 1021 1438 1023
rect 1446 1021 1449 1023
rect 1342 1012 1344 1021
rect 1432 1012 1434 1021
rect 816 1006 819 1008
rect 827 1006 837 1008
rect 730 1001 732 1004
rect 104 999 107 1001
rect 115 999 125 1001
rect 194 999 197 1001
rect 205 999 215 1001
rect 831 998 841 1000
rect 849 998 852 1000
rect -147 992 -137 994
rect -129 992 -126 994
rect -57 992 -47 994
rect -39 992 -36 994
rect -143 983 -141 992
rect -53 983 -51 992
rect 119 991 129 993
rect 137 991 140 993
rect 209 991 219 993
rect 227 991 230 993
rect 661 991 663 994
rect 691 992 693 995
rect 123 982 125 991
rect 213 982 215 991
rect 835 989 837 998
rect 1093 996 1106 998
rect 1114 996 1117 998
rect 1183 996 1196 998
rect 1204 996 1207 998
rect 1096 992 1098 996
rect 1186 992 1188 996
rect 1359 995 1372 997
rect 1380 995 1383 997
rect 1449 995 1462 997
rect 1470 995 1473 997
rect 1362 991 1364 995
rect 1452 991 1454 995
rect 661 979 663 983
rect 691 980 693 984
rect -182 971 -180 975
rect 661 977 672 979
rect -185 969 -172 971
rect -164 969 -161 971
rect 84 970 86 974
rect 661 973 663 977
rect 691 978 702 980
rect 691 974 693 978
rect 730 975 732 978
rect 81 968 94 970
rect 102 968 105 970
rect -126 966 -113 968
rect -105 966 -102 968
rect -36 966 -23 968
rect -15 966 -12 968
rect -123 962 -121 966
rect -205 953 -203 959
rect -33 962 -31 966
rect 140 965 153 967
rect 161 965 164 967
rect 230 965 243 967
rect 251 965 254 967
rect 653 968 655 971
rect 647 966 655 968
rect 852 972 865 974
rect 873 972 876 974
rect 855 968 857 972
rect 143 961 145 965
rect -221 951 -218 953
rect -210 951 -200 953
rect 61 952 63 958
rect 233 961 235 965
rect 653 961 655 966
rect 350 953 352 957
rect 730 959 732 967
rect 1046 967 1048 970
rect 722 957 732 959
rect 730 955 732 957
rect 45 950 48 952
rect 56 950 66 952
rect 347 951 360 953
rect 368 951 371 953
rect 623 950 625 953
rect 653 950 655 953
rect 402 945 404 948
rect -206 943 -196 945
rect -188 943 -185 945
rect -202 934 -200 943
rect 60 942 70 944
rect 78 942 81 944
rect 64 933 66 942
rect 327 935 329 941
rect 1046 951 1048 959
rect 1038 949 1048 951
rect 1046 947 1048 949
rect 730 944 732 947
rect 623 938 625 942
rect 311 933 314 935
rect 322 933 332 935
rect 326 925 336 927
rect 344 925 347 927
rect 402 929 404 937
rect 623 936 634 938
rect 623 932 625 936
rect 1046 936 1048 939
rect 394 927 404 929
rect 402 925 404 927
rect -185 917 -172 919
rect -164 917 -161 919
rect -182 913 -180 917
rect 81 916 94 918
rect 102 916 105 918
rect 330 916 332 925
rect 615 927 617 930
rect 609 925 617 927
rect 615 920 617 925
rect 84 912 86 916
rect 402 914 404 917
rect 730 918 732 921
rect 785 918 787 921
rect 1100 920 1102 924
rect 1190 920 1192 924
rect 1097 918 1110 920
rect 1118 918 1121 920
rect 1187 918 1200 920
rect 1208 918 1211 920
rect 1366 919 1368 923
rect 1456 919 1458 923
rect 585 909 587 912
rect 615 909 617 912
rect 1363 917 1376 919
rect 1384 917 1387 919
rect 1453 917 1466 919
rect 1474 917 1477 919
rect 347 899 360 901
rect 368 899 371 901
rect 350 895 352 899
rect 585 897 587 901
rect 730 902 732 910
rect 722 900 732 902
rect 730 898 732 900
rect 785 902 787 910
rect 1077 902 1079 908
rect 1167 902 1169 908
rect 777 900 787 902
rect 1061 900 1064 902
rect 1072 900 1082 902
rect 1151 900 1154 902
rect 1162 900 1172 902
rect 1343 901 1345 907
rect 1433 901 1435 907
rect 785 898 787 900
rect 1327 899 1330 901
rect 1338 899 1348 901
rect 1417 899 1420 901
rect 1428 899 1438 901
rect 585 895 596 897
rect 585 891 587 895
rect -127 878 -125 882
rect -37 878 -35 882
rect -130 876 -117 878
rect -109 876 -106 878
rect -40 876 -27 878
rect -19 876 -16 878
rect 139 877 141 881
rect 577 886 579 889
rect 730 887 732 890
rect 785 887 787 890
rect 855 888 857 892
rect 1076 892 1086 894
rect 1094 892 1097 894
rect 1166 892 1176 894
rect 1184 892 1187 894
rect 852 886 865 888
rect 873 886 876 888
rect 571 884 579 886
rect 229 877 231 881
rect 577 879 579 884
rect 1080 883 1082 892
rect 1170 883 1172 892
rect 1342 891 1352 893
rect 1360 891 1363 893
rect 1432 891 1442 893
rect 1450 891 1453 893
rect 136 875 149 877
rect 157 875 160 877
rect 226 875 239 877
rect 247 875 250 877
rect 547 875 549 878
rect 541 873 549 875
rect -150 860 -148 866
rect -60 860 -58 866
rect 547 868 549 873
rect 1346 882 1348 891
rect 1436 882 1438 891
rect 577 868 579 871
rect 832 870 834 876
rect 1041 871 1043 875
rect 816 868 819 870
rect 827 868 837 870
rect 1038 869 1051 871
rect 1059 869 1062 871
rect 1307 870 1309 874
rect 1304 868 1317 870
rect 1325 868 1328 870
rect -166 858 -163 860
rect -155 858 -145 860
rect -76 858 -73 860
rect -65 858 -55 860
rect 116 859 118 865
rect 206 859 208 865
rect 730 861 732 864
rect 1097 866 1110 868
rect 1118 866 1121 868
rect 1187 866 1200 868
rect 1208 866 1211 868
rect 100 857 103 859
rect 111 857 121 859
rect 190 857 193 859
rect 201 857 211 859
rect 325 856 327 859
rect 547 857 549 860
rect -151 850 -141 852
rect -133 850 -130 852
rect -61 850 -51 852
rect -43 850 -40 852
rect -147 841 -145 850
rect -57 841 -55 850
rect 115 849 125 851
rect 133 849 136 851
rect 205 849 215 851
rect 223 849 226 851
rect 119 840 121 849
rect 209 840 211 849
rect 831 860 841 862
rect 849 860 852 862
rect 325 840 327 848
rect 539 846 541 849
rect 533 844 541 846
rect 317 838 327 840
rect 539 839 541 844
rect 730 845 732 853
rect 835 851 837 860
rect 1100 862 1102 866
rect 1018 853 1020 859
rect 1190 862 1192 866
rect 1363 865 1376 867
rect 1384 865 1387 867
rect 1453 865 1466 867
rect 1474 865 1477 867
rect 1366 861 1368 865
rect 1002 851 1005 853
rect 1013 851 1023 853
rect 1284 852 1286 858
rect 1456 861 1458 865
rect 1268 850 1271 852
rect 1279 850 1289 852
rect 722 843 732 845
rect 941 843 943 847
rect 1017 843 1027 845
rect 1035 843 1038 845
rect 730 841 732 843
rect 938 841 951 843
rect 959 841 962 843
rect 325 836 327 838
rect -130 824 -117 826
rect -109 824 -106 826
rect -40 824 -27 826
rect -19 824 -16 826
rect 852 834 865 836
rect 873 834 876 836
rect 325 825 327 828
rect 395 826 397 830
rect 539 828 541 831
rect 730 830 732 833
rect 855 830 857 834
rect -127 820 -125 824
rect -37 820 -35 824
rect 136 823 149 825
rect 157 823 160 825
rect 226 823 239 825
rect 247 823 250 825
rect 392 824 405 826
rect 413 824 416 826
rect 1021 834 1023 843
rect 1283 842 1293 844
rect 1301 842 1304 844
rect 918 825 920 831
rect 1287 833 1289 842
rect 139 819 141 823
rect 229 819 231 823
rect 531 817 533 820
rect 525 815 533 817
rect 795 816 797 824
rect 902 823 905 825
rect 913 823 923 825
rect 1038 817 1051 819
rect 1059 817 1062 819
rect 372 808 374 814
rect 531 810 533 815
rect 782 814 785 816
rect 793 814 805 816
rect 813 814 816 816
rect 917 815 927 817
rect 935 815 938 817
rect 356 806 359 808
rect 367 806 377 808
rect 921 806 923 815
rect 1041 813 1043 817
rect 1304 816 1317 818
rect 1325 816 1328 818
rect 1307 812 1309 816
rect 371 798 381 800
rect 389 798 392 800
rect 531 799 533 802
rect -177 795 -175 798
rect 375 789 377 798
rect 855 793 857 797
rect 852 791 865 793
rect 873 791 876 793
rect -177 779 -175 787
rect 938 789 951 791
rect 959 789 962 791
rect 481 781 483 785
rect 941 785 943 789
rect 478 779 491 781
rect 499 779 502 781
rect -185 777 -175 779
rect -177 775 -175 777
rect 832 775 834 781
rect 1096 778 1098 782
rect 1186 778 1188 782
rect 1093 776 1106 778
rect 1114 776 1117 778
rect 1183 776 1196 778
rect 1204 776 1207 778
rect 1362 777 1364 781
rect 1452 777 1454 781
rect 392 772 405 774
rect 413 772 416 774
rect 816 773 819 775
rect 827 773 837 775
rect 395 768 397 772
rect -177 764 -175 767
rect 458 763 460 769
rect 1359 775 1372 777
rect 1380 775 1383 777
rect 1449 775 1462 777
rect 1470 775 1473 777
rect 831 765 841 767
rect 849 765 852 767
rect -123 748 -121 752
rect -33 748 -31 752
rect -126 746 -113 748
rect -105 746 -102 748
rect -36 746 -23 748
rect -15 746 -12 748
rect 143 747 145 751
rect 335 754 337 762
rect 442 761 445 763
rect 453 761 463 763
rect 835 756 837 765
rect 1073 760 1075 766
rect 1163 760 1165 766
rect 1057 758 1060 760
rect 1068 758 1078 760
rect 1147 758 1150 760
rect 1158 758 1168 760
rect 1339 759 1341 765
rect 1429 759 1431 765
rect 1323 757 1326 759
rect 1334 757 1344 759
rect 1413 757 1416 759
rect 1424 757 1434 759
rect 322 752 325 754
rect 333 752 345 754
rect 353 752 356 754
rect 457 753 467 755
rect 475 753 478 755
rect 233 747 235 751
rect 140 745 153 747
rect 161 745 164 747
rect 230 745 243 747
rect 251 745 254 747
rect 461 744 463 753
rect 1072 750 1082 752
rect 1090 750 1093 752
rect 1162 750 1172 752
rect 1180 750 1183 752
rect 1076 741 1078 750
rect 1166 741 1168 750
rect 1338 749 1348 751
rect 1356 749 1359 751
rect 1428 749 1438 751
rect 1446 749 1449 751
rect 852 739 865 741
rect 873 739 876 741
rect -146 730 -144 736
rect -56 730 -54 736
rect -162 728 -159 730
rect -151 728 -141 730
rect -72 728 -69 730
rect -61 728 -51 730
rect 120 729 122 735
rect 210 729 212 735
rect 395 731 397 735
rect 855 735 857 739
rect 392 729 405 731
rect 413 729 416 731
rect 1342 740 1344 749
rect 1432 740 1434 749
rect 104 727 107 729
rect 115 727 125 729
rect 194 727 197 729
rect 205 727 215 729
rect 478 727 491 729
rect 499 727 502 729
rect 481 723 483 727
rect -147 720 -137 722
rect -129 720 -126 722
rect -57 720 -47 722
rect -39 720 -36 722
rect -143 711 -141 720
rect -53 711 -51 720
rect 119 719 129 721
rect 137 719 140 721
rect 209 719 219 721
rect 227 719 230 721
rect 1093 724 1106 726
rect 1114 724 1117 726
rect 1183 724 1196 726
rect 1204 724 1207 726
rect 1096 720 1098 724
rect 123 710 125 719
rect 213 710 215 719
rect 372 713 374 719
rect 1186 720 1188 724
rect 1359 723 1372 725
rect 1380 723 1383 725
rect 1449 723 1462 725
rect 1470 723 1473 725
rect 1362 719 1364 723
rect 1452 719 1454 723
rect 356 711 359 713
rect 367 711 377 713
rect -182 699 -180 703
rect 371 703 381 705
rect 389 703 392 705
rect -185 697 -172 699
rect -164 697 -161 699
rect 84 698 86 702
rect 81 696 94 698
rect 102 696 105 698
rect -126 694 -113 696
rect -105 694 -102 696
rect -36 694 -23 696
rect -15 694 -12 696
rect -123 690 -121 694
rect -205 681 -203 687
rect -33 690 -31 694
rect 140 693 153 695
rect 161 693 164 695
rect 230 693 243 695
rect 251 693 254 695
rect 375 694 377 703
rect 1046 695 1048 698
rect 143 689 145 693
rect -221 679 -218 681
rect -210 679 -200 681
rect 61 680 63 686
rect 233 689 235 693
rect 785 685 787 688
rect 45 678 48 680
rect 56 678 66 680
rect 392 677 405 679
rect 413 677 416 679
rect 395 673 397 677
rect -206 671 -196 673
rect -188 671 -185 673
rect -202 662 -200 671
rect 60 670 70 672
rect 78 670 81 672
rect 64 661 66 670
rect 785 669 787 677
rect 1046 679 1048 687
rect 1038 677 1048 679
rect 1046 675 1048 677
rect 777 667 787 669
rect 785 665 787 667
rect 1046 664 1048 667
rect 785 654 787 657
rect 855 655 857 659
rect 852 653 865 655
rect 873 653 876 655
rect 1100 648 1102 652
rect 1190 648 1192 652
rect -185 645 -172 647
rect -164 645 -161 647
rect -182 641 -180 645
rect 81 644 94 646
rect 102 644 105 646
rect 84 640 86 644
rect 1097 646 1110 648
rect 1118 646 1121 648
rect 1187 646 1200 648
rect 1208 646 1211 648
rect 1366 647 1368 651
rect 1456 647 1458 651
rect 832 637 834 643
rect 1363 645 1376 647
rect 1384 645 1387 647
rect 1453 645 1466 647
rect 1474 645 1477 647
rect 816 635 819 637
rect 827 635 837 637
rect 1077 630 1079 636
rect 1167 630 1169 636
rect 831 627 841 629
rect 849 627 852 629
rect 1061 628 1064 630
rect 1072 628 1082 630
rect 1151 628 1154 630
rect 1162 628 1172 630
rect 1343 629 1345 635
rect 1433 629 1435 635
rect 1327 627 1330 629
rect 1338 627 1348 629
rect 1417 627 1420 629
rect 1428 627 1438 629
rect 350 618 352 622
rect 835 618 837 627
rect 1076 620 1086 622
rect 1094 620 1097 622
rect 1166 620 1176 622
rect 1184 620 1187 622
rect 347 616 360 618
rect 368 616 371 618
rect -127 606 -125 610
rect -37 606 -35 610
rect -130 604 -117 606
rect -109 604 -106 606
rect -40 604 -27 606
rect -19 604 -16 606
rect 139 605 141 609
rect 402 610 404 613
rect 941 610 943 614
rect 1080 611 1082 620
rect 1170 611 1172 620
rect 1342 619 1352 621
rect 1360 619 1363 621
rect 1432 619 1442 621
rect 1450 619 1453 621
rect 229 605 231 609
rect 136 603 149 605
rect 157 603 160 605
rect 226 603 239 605
rect 247 603 250 605
rect 327 600 329 606
rect 938 608 951 610
rect 959 608 962 610
rect 1346 610 1348 619
rect 1436 610 1438 619
rect 311 598 314 600
rect 322 598 332 600
rect -150 588 -148 594
rect -60 588 -58 594
rect -166 586 -163 588
rect -155 586 -145 588
rect -76 586 -73 588
rect -65 586 -55 588
rect 116 587 118 593
rect 206 587 208 593
rect 326 590 336 592
rect 344 590 347 592
rect 402 594 404 602
rect 852 601 865 603
rect 873 601 876 603
rect 855 597 857 601
rect 394 592 404 594
rect 402 590 404 592
rect 1041 599 1043 603
rect 918 592 920 598
rect 1038 597 1051 599
rect 1059 597 1062 599
rect 1307 598 1309 602
rect 1304 596 1317 598
rect 1325 596 1328 598
rect 1097 594 1110 596
rect 1118 594 1121 596
rect 1187 594 1200 596
rect 1208 594 1211 596
rect 100 585 103 587
rect 111 585 121 587
rect 190 585 193 587
rect 201 585 211 587
rect 330 581 332 590
rect 795 583 797 591
rect 902 590 905 592
rect 913 590 923 592
rect 1100 590 1102 594
rect -151 578 -141 580
rect -133 578 -130 580
rect -61 578 -51 580
rect -43 578 -40 580
rect -147 569 -145 578
rect -57 569 -55 578
rect 115 577 125 579
rect 133 577 136 579
rect 205 577 215 579
rect 223 577 226 579
rect 402 579 404 582
rect 782 581 785 583
rect 793 581 805 583
rect 813 581 816 583
rect 917 582 927 584
rect 935 582 938 584
rect 119 568 121 577
rect 209 568 211 577
rect 921 573 923 582
rect 1018 581 1020 587
rect 1190 590 1192 594
rect 1363 593 1376 595
rect 1384 593 1387 595
rect 1453 593 1466 595
rect 1474 593 1477 595
rect 1366 589 1368 593
rect 1002 579 1005 581
rect 1013 579 1023 581
rect 1284 580 1286 586
rect 1456 589 1458 593
rect 1268 578 1271 580
rect 1279 578 1289 580
rect 1017 571 1027 573
rect 1035 571 1038 573
rect 347 564 360 566
rect 368 564 371 566
rect 350 560 352 564
rect -130 552 -117 554
rect -109 552 -106 554
rect -40 552 -27 554
rect -19 552 -16 554
rect 855 560 857 564
rect 852 558 865 560
rect 873 558 876 560
rect 1021 562 1023 571
rect 1283 570 1293 572
rect 1301 570 1304 572
rect 1287 561 1289 570
rect 938 556 951 558
rect 959 556 962 558
rect -127 548 -125 552
rect -37 548 -35 552
rect 136 551 149 553
rect 157 551 160 553
rect 226 551 239 553
rect 247 551 250 553
rect 941 552 943 556
rect 139 547 141 551
rect 229 547 231 551
rect 832 542 834 548
rect 1038 545 1051 547
rect 1059 545 1062 547
rect 816 540 819 542
rect 827 540 837 542
rect 1041 541 1043 545
rect 1304 544 1317 546
rect 1325 544 1328 546
rect 1307 540 1309 544
rect 831 532 841 534
rect 849 532 852 534
rect -177 523 -175 526
rect 325 521 327 524
rect 835 523 837 532
rect -177 507 -175 515
rect -185 505 -175 507
rect -177 503 -175 505
rect 325 505 327 513
rect 852 506 865 508
rect 873 506 876 508
rect 1096 506 1098 510
rect 1186 506 1188 510
rect 317 503 327 505
rect 325 501 327 503
rect 855 502 857 506
rect -177 492 -175 495
rect 1093 504 1106 506
rect 1114 504 1117 506
rect 1183 504 1196 506
rect 1204 504 1207 506
rect 1362 505 1364 509
rect 1452 505 1454 509
rect 1359 503 1372 505
rect 1380 503 1383 505
rect 1449 503 1462 505
rect 1470 503 1473 505
rect 325 490 327 493
rect 395 491 397 495
rect 392 489 405 491
rect 413 489 416 491
rect 1073 488 1075 494
rect 1163 488 1165 494
rect 1057 486 1060 488
rect 1068 486 1078 488
rect 1147 486 1150 488
rect 1158 486 1168 488
rect 1339 487 1341 493
rect 1429 487 1431 493
rect 1323 485 1326 487
rect 1334 485 1344 487
rect 1413 485 1416 487
rect 1424 485 1434 487
rect -123 476 -121 480
rect -33 476 -31 480
rect -126 474 -113 476
rect -105 474 -102 476
rect -36 474 -23 476
rect -15 474 -12 476
rect 143 475 145 479
rect 233 475 235 479
rect 140 473 153 475
rect 161 473 164 475
rect 230 473 243 475
rect 251 473 254 475
rect 372 473 374 479
rect 1072 478 1082 480
rect 1090 478 1093 480
rect 1162 478 1172 480
rect 1180 478 1183 480
rect 356 471 359 473
rect 367 471 377 473
rect -146 458 -144 464
rect -56 458 -54 464
rect 1076 469 1078 478
rect 1166 469 1168 478
rect 1338 477 1348 479
rect 1356 477 1359 479
rect 1428 477 1438 479
rect 1446 477 1449 479
rect 1342 468 1344 477
rect 1432 468 1434 477
rect 371 463 381 465
rect 389 463 392 465
rect -162 456 -159 458
rect -151 456 -141 458
rect -72 456 -69 458
rect -61 456 -51 458
rect 120 457 122 463
rect 210 457 212 463
rect 104 455 107 457
rect 115 455 125 457
rect 194 455 197 457
rect 205 455 215 457
rect 375 454 377 463
rect 1093 452 1106 454
rect 1114 452 1117 454
rect 1183 452 1196 454
rect 1204 452 1207 454
rect -147 448 -137 450
rect -129 448 -126 450
rect -57 448 -47 450
rect -39 448 -36 450
rect -143 439 -141 448
rect -53 439 -51 448
rect 119 447 129 449
rect 137 447 140 449
rect 209 447 219 449
rect 227 447 230 449
rect 123 438 125 447
rect 213 438 215 447
rect 481 446 483 450
rect 1096 448 1098 452
rect 478 444 491 446
rect 499 444 502 446
rect 1186 448 1188 452
rect 1359 451 1372 453
rect 1380 451 1383 453
rect 1449 451 1462 453
rect 1470 451 1473 453
rect 1362 447 1364 451
rect 1452 447 1454 451
rect 392 437 405 439
rect 413 437 416 439
rect -182 427 -180 431
rect 395 433 397 437
rect -185 425 -172 427
rect -164 425 -161 427
rect 84 426 86 430
rect 81 424 94 426
rect 102 424 105 426
rect -126 422 -113 424
rect -105 422 -102 424
rect -36 422 -23 424
rect -15 422 -12 424
rect 458 428 460 434
rect -123 418 -121 422
rect -205 409 -203 415
rect -33 418 -31 422
rect 140 421 153 423
rect 161 421 164 423
rect 230 421 243 423
rect 251 421 254 423
rect 143 417 145 421
rect -221 407 -218 409
rect -210 407 -200 409
rect 61 408 63 414
rect 233 417 235 421
rect 335 419 337 427
rect 442 426 445 428
rect 453 426 463 428
rect 1046 423 1048 426
rect 322 417 325 419
rect 333 417 345 419
rect 353 417 356 419
rect 457 418 467 420
rect 475 418 478 420
rect 461 409 463 418
rect 45 406 48 408
rect 56 406 66 408
rect 1046 407 1048 415
rect 1038 405 1048 407
rect -206 399 -196 401
rect -188 399 -185 401
rect 1046 403 1048 405
rect -202 390 -200 399
rect 60 398 70 400
rect 78 398 81 400
rect 64 389 66 398
rect 395 396 397 400
rect 392 394 405 396
rect 413 394 416 396
rect 478 392 491 394
rect 499 392 502 394
rect 1046 392 1048 395
rect 481 388 483 392
rect 372 378 374 384
rect 356 376 359 378
rect 367 376 377 378
rect 1100 376 1102 380
rect 1190 376 1192 380
rect -185 373 -172 375
rect -164 373 -161 375
rect -182 369 -180 373
rect 81 372 94 374
rect 102 372 105 374
rect 84 368 86 372
rect 1097 374 1110 376
rect 1118 374 1121 376
rect 1187 374 1200 376
rect 1208 374 1211 376
rect 1366 375 1368 379
rect 1456 375 1458 379
rect 371 368 381 370
rect 389 368 392 370
rect 1363 373 1376 375
rect 1384 373 1387 375
rect 1453 373 1466 375
rect 1474 373 1477 375
rect 375 359 377 368
rect 1077 358 1079 364
rect 1167 358 1169 364
rect 1061 356 1064 358
rect 1072 356 1082 358
rect 1151 356 1154 358
rect 1162 356 1172 358
rect 1343 357 1345 363
rect 1433 357 1435 363
rect 1327 355 1330 357
rect 1338 355 1348 357
rect 1417 355 1420 357
rect 1428 355 1438 357
rect 1076 348 1086 350
rect 1094 348 1097 350
rect 1166 348 1176 350
rect 1184 348 1187 350
rect 392 342 405 344
rect 413 342 416 344
rect -127 334 -125 338
rect -37 334 -35 338
rect -130 332 -117 334
rect -109 332 -106 334
rect -40 332 -27 334
rect -19 332 -16 334
rect 139 333 141 337
rect 395 338 397 342
rect 229 333 231 337
rect 1080 339 1082 348
rect 1170 339 1172 348
rect 1342 347 1352 349
rect 1360 347 1363 349
rect 1432 347 1442 349
rect 1450 347 1453 349
rect 1346 338 1348 347
rect 1436 338 1438 347
rect 136 331 149 333
rect 157 331 160 333
rect 226 331 239 333
rect 247 331 250 333
rect 1041 327 1043 331
rect 1038 325 1051 327
rect 1059 325 1062 327
rect -150 316 -148 322
rect -60 316 -58 322
rect 1307 326 1309 330
rect 1304 324 1317 326
rect 1325 324 1328 326
rect -166 314 -163 316
rect -155 314 -145 316
rect -76 314 -73 316
rect -65 314 -55 316
rect 116 315 118 321
rect 206 315 208 321
rect 1097 322 1110 324
rect 1118 322 1121 324
rect 1187 322 1200 324
rect 1208 322 1211 324
rect 1100 318 1102 322
rect 100 313 103 315
rect 111 313 121 315
rect 190 313 193 315
rect 201 313 211 315
rect 1018 309 1020 315
rect 1190 318 1192 322
rect 1363 321 1376 323
rect 1384 321 1387 323
rect 1453 321 1466 323
rect 1474 321 1477 323
rect 1366 317 1368 321
rect -151 306 -141 308
rect -133 306 -130 308
rect -61 306 -51 308
rect -43 306 -40 308
rect 1002 307 1005 309
rect 1013 307 1023 309
rect 1284 308 1286 314
rect 1456 317 1458 321
rect -147 297 -145 306
rect -57 297 -55 306
rect 115 305 125 307
rect 133 305 136 307
rect 205 305 215 307
rect 223 305 226 307
rect 1268 306 1271 308
rect 1279 306 1289 308
rect 119 296 121 305
rect 209 296 211 305
rect 1017 299 1027 301
rect 1035 299 1038 301
rect 1021 290 1023 299
rect 1283 298 1293 300
rect 1301 298 1304 300
rect -130 280 -117 282
rect -109 280 -106 282
rect -40 280 -27 282
rect -19 280 -16 282
rect 350 283 352 287
rect 1287 289 1289 298
rect 347 281 360 283
rect 368 281 371 283
rect -127 276 -125 280
rect -37 276 -35 280
rect 136 279 149 281
rect 157 279 160 281
rect 226 279 239 281
rect 247 279 250 281
rect 139 275 141 279
rect 229 275 231 279
rect 402 275 404 278
rect 327 265 329 271
rect 1038 273 1051 275
rect 1059 273 1062 275
rect 1041 269 1043 273
rect 1304 272 1317 274
rect 1325 272 1328 274
rect 311 263 314 265
rect 322 263 332 265
rect 326 255 336 257
rect 344 255 347 257
rect 402 259 404 267
rect 1307 268 1309 272
rect 394 257 404 259
rect 402 255 404 257
rect -177 251 -175 254
rect 330 246 332 255
rect -177 235 -175 243
rect 402 244 404 247
rect -185 233 -175 235
rect -177 231 -175 233
rect 347 229 360 231
rect 368 229 371 231
rect 350 225 352 229
rect -177 220 -175 223
rect -123 204 -121 208
rect -33 204 -31 208
rect -126 202 -113 204
rect -105 202 -102 204
rect -36 202 -23 204
rect -15 202 -12 204
rect 143 203 145 207
rect 233 203 235 207
rect 140 201 153 203
rect 161 201 164 203
rect 230 201 243 203
rect 251 201 254 203
rect -146 186 -144 192
rect -56 186 -54 192
rect -162 184 -159 186
rect -151 184 -141 186
rect -72 184 -69 186
rect -61 184 -51 186
rect 120 185 122 191
rect 210 185 212 191
rect 104 183 107 185
rect 115 183 125 185
rect 194 183 197 185
rect 205 183 215 185
rect -147 176 -137 178
rect -129 176 -126 178
rect -57 176 -47 178
rect -39 176 -36 178
rect -143 167 -141 176
rect -53 167 -51 176
rect 119 175 129 177
rect 137 175 140 177
rect 209 175 219 177
rect 227 175 230 177
rect 123 166 125 175
rect 213 166 215 175
rect -182 155 -180 159
rect -185 153 -172 155
rect -164 153 -161 155
rect 84 154 86 158
rect 81 152 94 154
rect 102 152 105 154
rect -126 150 -113 152
rect -105 150 -102 152
rect -36 150 -23 152
rect -15 150 -12 152
rect -123 146 -121 150
rect -205 137 -203 143
rect -33 146 -31 150
rect 140 149 153 151
rect 161 149 164 151
rect 230 149 243 151
rect 251 149 254 151
rect 143 145 145 149
rect -221 135 -218 137
rect -210 135 -200 137
rect 61 136 63 142
rect 233 145 235 149
rect 45 134 48 136
rect 56 134 66 136
rect -206 127 -196 129
rect -188 127 -185 129
rect -202 118 -200 127
rect 60 126 70 128
rect 78 126 81 128
rect 64 117 66 126
rect -185 101 -172 103
rect -164 101 -161 103
rect -182 97 -180 101
rect 81 100 94 102
rect 102 100 105 102
rect 84 96 86 100
rect -127 62 -125 66
rect -37 62 -35 66
rect -130 60 -117 62
rect -109 60 -106 62
rect -40 60 -27 62
rect -19 60 -16 62
rect 139 61 141 65
rect 229 61 231 65
rect 136 59 149 61
rect 157 59 160 61
rect 226 59 239 61
rect 247 59 250 61
rect -150 44 -148 50
rect -60 44 -58 50
rect -166 42 -163 44
rect -155 42 -145 44
rect -76 42 -73 44
rect -65 42 -55 44
rect 116 43 118 49
rect 206 43 208 49
rect 100 41 103 43
rect 111 41 121 43
rect 190 41 193 43
rect 201 41 211 43
rect -151 34 -141 36
rect -133 34 -130 36
rect -61 34 -51 36
rect -43 34 -40 36
rect -147 25 -145 34
rect -57 25 -55 34
rect 115 33 125 35
rect 133 33 136 35
rect 205 33 215 35
rect 223 33 226 35
rect 119 24 121 33
rect 209 24 211 33
rect -130 8 -117 10
rect -109 8 -106 10
rect -40 8 -27 10
rect -19 8 -16 10
rect -127 4 -125 8
rect -37 4 -35 8
rect 136 7 149 9
rect 157 7 160 9
rect 226 7 239 9
rect 247 7 250 9
rect 139 3 141 7
rect 229 3 231 7
rect -177 -21 -175 -18
rect -177 -37 -175 -29
rect -185 -39 -175 -37
rect -177 -41 -175 -39
rect -177 -52 -175 -49
rect -123 -68 -121 -64
rect -33 -68 -31 -64
rect -126 -70 -113 -68
rect -105 -70 -102 -68
rect -36 -70 -23 -68
rect -15 -70 -12 -68
rect 143 -69 145 -65
rect 233 -69 235 -65
rect 140 -71 153 -69
rect 161 -71 164 -69
rect 230 -71 243 -69
rect 251 -71 254 -69
rect -146 -86 -144 -80
rect -56 -86 -54 -80
rect -162 -88 -159 -86
rect -151 -88 -141 -86
rect -72 -88 -69 -86
rect -61 -88 -51 -86
rect 120 -87 122 -81
rect 210 -87 212 -81
rect 104 -89 107 -87
rect 115 -89 125 -87
rect 194 -89 197 -87
rect 205 -89 215 -87
rect -147 -96 -137 -94
rect -129 -96 -126 -94
rect -57 -96 -47 -94
rect -39 -96 -36 -94
rect -143 -105 -141 -96
rect -53 -105 -51 -96
rect 119 -97 129 -95
rect 137 -97 140 -95
rect 209 -97 219 -95
rect 227 -97 230 -95
rect 123 -106 125 -97
rect 213 -106 215 -97
rect -182 -117 -180 -113
rect -185 -119 -172 -117
rect -164 -119 -161 -117
rect 84 -118 86 -114
rect 81 -120 94 -118
rect 102 -120 105 -118
rect -126 -122 -113 -120
rect -105 -122 -102 -120
rect -36 -122 -23 -120
rect -15 -122 -12 -120
rect -123 -126 -121 -122
rect -205 -135 -203 -129
rect -33 -126 -31 -122
rect 140 -123 153 -121
rect 161 -123 164 -121
rect 230 -123 243 -121
rect 251 -123 254 -121
rect 143 -127 145 -123
rect -221 -137 -218 -135
rect -210 -137 -200 -135
rect 61 -136 63 -130
rect 233 -127 235 -123
rect 45 -138 48 -136
rect 56 -138 66 -136
rect -206 -145 -196 -143
rect -188 -145 -185 -143
rect -202 -154 -200 -145
rect 60 -146 70 -144
rect 78 -146 81 -144
rect 64 -155 66 -146
rect -185 -171 -172 -169
rect -164 -171 -161 -169
rect -182 -175 -180 -171
rect 81 -172 94 -170
rect 102 -172 105 -170
rect 84 -176 86 -172
<< polycontact >>
rect -128 1970 -124 1974
rect -38 1970 -34 1974
rect 138 1969 142 1973
rect 228 1969 232 1973
rect -151 1954 -147 1958
rect -61 1954 -57 1958
rect 115 1953 119 1957
rect 205 1953 209 1957
rect -148 1925 -144 1929
rect -58 1925 -54 1929
rect 118 1924 122 1928
rect 208 1924 212 1928
rect -128 1904 -124 1908
rect -38 1904 -34 1908
rect 138 1903 142 1907
rect 228 1903 232 1907
rect -189 1864 -185 1868
rect -124 1840 -120 1844
rect -34 1840 -30 1844
rect 142 1839 146 1843
rect 232 1839 236 1843
rect -147 1824 -143 1828
rect -57 1824 -53 1828
rect 119 1823 123 1827
rect 209 1823 213 1827
rect -144 1795 -140 1799
rect -54 1795 -50 1799
rect -183 1791 -179 1795
rect 122 1794 126 1798
rect 212 1794 216 1798
rect 83 1790 87 1794
rect -206 1775 -202 1779
rect -124 1774 -120 1778
rect -34 1774 -30 1778
rect 60 1774 64 1778
rect 142 1773 146 1777
rect 232 1773 236 1777
rect -203 1746 -199 1750
rect 63 1745 67 1749
rect -183 1725 -179 1729
rect 83 1724 87 1728
rect -128 1698 -124 1702
rect -38 1698 -34 1702
rect 138 1697 142 1701
rect 228 1697 232 1701
rect -151 1682 -147 1686
rect -61 1682 -57 1686
rect 115 1681 119 1685
rect 205 1681 209 1685
rect -148 1653 -144 1657
rect -58 1653 -54 1657
rect 118 1652 122 1656
rect 208 1652 212 1656
rect -128 1632 -124 1636
rect -38 1632 -34 1636
rect 138 1631 142 1635
rect 228 1631 232 1635
rect -189 1592 -185 1596
rect 1095 1598 1099 1602
rect 1185 1598 1189 1602
rect 1361 1597 1365 1601
rect 1451 1597 1455 1601
rect 1072 1582 1076 1586
rect 1162 1582 1166 1586
rect 1338 1581 1342 1585
rect 1428 1581 1432 1585
rect -124 1568 -120 1572
rect -34 1568 -30 1572
rect 142 1567 146 1571
rect 232 1567 236 1571
rect -147 1552 -143 1556
rect -57 1552 -53 1556
rect 119 1551 123 1555
rect 209 1551 213 1555
rect 1075 1553 1079 1557
rect 1165 1553 1169 1557
rect 1341 1552 1345 1556
rect 1431 1552 1435 1556
rect -144 1523 -140 1527
rect -54 1523 -50 1527
rect 1095 1532 1099 1536
rect 1185 1532 1189 1536
rect 1361 1531 1365 1535
rect 1451 1531 1455 1535
rect -183 1519 -179 1523
rect 122 1522 126 1526
rect 212 1522 216 1526
rect 83 1518 87 1522
rect -206 1503 -202 1507
rect -124 1502 -120 1506
rect -34 1502 -30 1506
rect 60 1502 64 1506
rect 142 1501 146 1505
rect 232 1501 236 1505
rect 313 1507 317 1511
rect 394 1500 398 1504
rect 1034 1492 1038 1496
rect -203 1474 -199 1478
rect 371 1484 375 1488
rect 63 1473 67 1477
rect 1099 1468 1103 1472
rect -183 1453 -179 1457
rect 1189 1468 1193 1472
rect 1365 1467 1369 1471
rect 1455 1467 1459 1471
rect 83 1452 87 1456
rect 374 1455 378 1459
rect 480 1455 484 1459
rect 1076 1452 1080 1456
rect 1166 1452 1170 1456
rect 1342 1451 1346 1455
rect 1432 1451 1436 1455
rect 334 1432 338 1436
rect 394 1434 398 1438
rect 457 1439 461 1443
rect -128 1426 -124 1430
rect -38 1426 -34 1430
rect 138 1425 142 1429
rect 228 1425 232 1429
rect 1079 1423 1083 1427
rect 1169 1423 1173 1427
rect 1040 1419 1044 1423
rect 1345 1422 1349 1426
rect 1435 1422 1439 1426
rect 1306 1418 1310 1422
rect -151 1410 -147 1414
rect -61 1410 -57 1414
rect 115 1409 119 1413
rect 205 1409 209 1413
rect 460 1410 464 1414
rect 394 1405 398 1409
rect 1017 1403 1021 1407
rect 1099 1402 1103 1406
rect 1189 1402 1193 1406
rect 1283 1402 1287 1406
rect -148 1381 -144 1385
rect -58 1381 -54 1385
rect 371 1389 375 1393
rect 480 1389 484 1393
rect 1365 1401 1369 1405
rect 1455 1401 1459 1405
rect 118 1380 122 1384
rect 208 1380 212 1384
rect -128 1360 -124 1364
rect -38 1360 -34 1364
rect 138 1359 142 1363
rect 228 1359 232 1363
rect 773 1365 777 1369
rect 1020 1374 1024 1378
rect 1286 1373 1290 1377
rect 374 1360 378 1364
rect 854 1358 858 1362
rect 1040 1353 1044 1357
rect 1306 1352 1310 1356
rect 394 1339 398 1343
rect 831 1342 835 1346
rect -189 1320 -185 1324
rect 1095 1326 1099 1330
rect 1185 1326 1189 1330
rect 1361 1325 1365 1329
rect 1451 1325 1455 1329
rect 834 1313 838 1317
rect 940 1313 944 1317
rect 1072 1310 1076 1314
rect 1162 1310 1166 1314
rect 1338 1309 1342 1313
rect 1428 1309 1432 1313
rect -124 1296 -120 1300
rect -34 1296 -30 1300
rect 142 1295 146 1299
rect 232 1295 236 1299
rect 349 1292 353 1296
rect 794 1290 798 1294
rect 854 1292 858 1296
rect 917 1297 921 1301
rect -147 1280 -143 1284
rect -57 1280 -53 1284
rect 119 1279 123 1283
rect 209 1279 213 1283
rect 1075 1281 1079 1285
rect 1165 1281 1169 1285
rect 326 1276 330 1280
rect 1341 1280 1345 1284
rect 1431 1280 1435 1284
rect -144 1251 -140 1255
rect -54 1251 -50 1255
rect 390 1261 394 1265
rect 920 1268 924 1272
rect 854 1263 858 1267
rect -183 1247 -179 1251
rect 122 1250 126 1254
rect 212 1250 216 1254
rect 1095 1260 1099 1264
rect 1185 1260 1189 1264
rect 1361 1259 1365 1263
rect 1451 1259 1455 1263
rect 83 1246 87 1250
rect 329 1247 333 1251
rect 831 1247 835 1251
rect 940 1247 944 1251
rect -206 1231 -202 1235
rect -124 1230 -120 1234
rect -34 1230 -30 1234
rect 60 1230 64 1234
rect 142 1229 146 1233
rect 232 1229 236 1233
rect 349 1226 353 1230
rect 834 1218 838 1222
rect 1034 1220 1038 1224
rect -203 1202 -199 1206
rect 63 1201 67 1205
rect 854 1197 858 1201
rect 1099 1196 1103 1200
rect 1189 1196 1193 1200
rect 1365 1195 1369 1199
rect -183 1181 -179 1185
rect 83 1180 87 1184
rect 1455 1195 1459 1199
rect 313 1172 317 1176
rect 1076 1180 1080 1184
rect 1166 1180 1170 1184
rect 1342 1179 1346 1183
rect 1432 1179 1436 1183
rect 394 1165 398 1169
rect -128 1154 -124 1158
rect -38 1154 -34 1158
rect 138 1153 142 1157
rect 228 1153 232 1157
rect 371 1149 375 1153
rect 1079 1151 1083 1155
rect 1169 1151 1173 1155
rect 1040 1147 1044 1151
rect 1345 1150 1349 1154
rect 1435 1150 1439 1154
rect 1306 1146 1310 1150
rect -151 1138 -147 1142
rect -61 1138 -57 1142
rect 115 1137 119 1141
rect 205 1137 209 1141
rect 773 1132 777 1136
rect 1017 1131 1021 1135
rect -148 1109 -144 1113
rect -58 1109 -54 1113
rect 374 1120 378 1124
rect 480 1120 484 1124
rect 854 1125 858 1129
rect 1099 1130 1103 1134
rect 1189 1130 1193 1134
rect 1283 1130 1287 1134
rect 1365 1129 1369 1133
rect 1455 1129 1459 1133
rect 118 1108 122 1112
rect 208 1108 212 1112
rect 831 1109 835 1113
rect 334 1097 338 1101
rect 394 1099 398 1103
rect 457 1104 461 1108
rect 1020 1102 1024 1106
rect 1286 1101 1290 1105
rect -128 1088 -124 1092
rect -38 1088 -34 1092
rect 138 1087 142 1091
rect 228 1087 232 1091
rect 834 1080 838 1084
rect 940 1080 944 1084
rect 1040 1081 1044 1085
rect 460 1075 464 1079
rect 1306 1080 1310 1084
rect 394 1070 398 1074
rect -189 1048 -185 1052
rect 371 1054 375 1058
rect 480 1054 484 1058
rect 794 1057 798 1061
rect 854 1059 858 1063
rect 917 1064 921 1068
rect 1095 1054 1099 1058
rect 1185 1054 1189 1058
rect 1361 1053 1365 1057
rect 1451 1053 1455 1057
rect 920 1035 924 1039
rect 1072 1038 1076 1042
rect 1162 1038 1166 1042
rect -124 1024 -120 1028
rect -34 1024 -30 1028
rect 142 1023 146 1027
rect 232 1023 236 1027
rect 374 1025 378 1029
rect 854 1030 858 1034
rect 1338 1037 1342 1041
rect 1428 1037 1432 1041
rect 539 1012 543 1016
rect -147 1008 -143 1012
rect -57 1008 -53 1012
rect 119 1007 123 1011
rect 209 1007 213 1011
rect 394 1004 398 1008
rect 577 1012 581 1016
rect 615 1012 619 1016
rect 653 1012 657 1016
rect 718 1013 722 1017
rect 831 1014 835 1018
rect 940 1014 944 1018
rect 1075 1009 1079 1013
rect 1165 1009 1169 1013
rect 1341 1008 1345 1012
rect 1431 1008 1435 1012
rect -144 979 -140 983
rect -54 979 -50 983
rect 834 985 838 989
rect 1095 988 1099 992
rect 1185 988 1189 992
rect 1361 987 1365 991
rect 1451 987 1455 991
rect -183 975 -179 979
rect 122 978 126 982
rect 212 978 216 982
rect 83 974 87 978
rect 672 976 676 980
rect 702 977 706 981
rect -206 959 -202 963
rect -124 958 -120 962
rect -34 958 -30 962
rect 643 965 647 969
rect 60 958 64 962
rect 142 957 146 961
rect 232 957 236 961
rect 349 957 353 961
rect 718 956 722 960
rect 854 964 858 968
rect -203 930 -199 934
rect 326 941 330 945
rect 1034 948 1038 952
rect 63 929 67 933
rect 390 926 394 930
rect 634 935 638 939
rect 605 924 609 928
rect 1099 924 1103 928
rect -183 909 -179 913
rect 83 908 87 912
rect 329 912 333 916
rect 1189 924 1193 928
rect 1365 923 1369 927
rect 1455 923 1459 927
rect 349 891 353 895
rect 718 899 722 903
rect 773 899 777 903
rect 1076 908 1080 912
rect 1166 908 1170 912
rect 1342 907 1346 911
rect 1432 907 1436 911
rect 596 894 600 898
rect 854 892 858 896
rect -128 882 -124 886
rect -38 882 -34 886
rect 138 881 142 885
rect 228 881 232 885
rect 567 883 571 887
rect 537 872 541 876
rect -151 866 -147 870
rect -61 866 -57 870
rect 115 865 119 869
rect 205 865 209 869
rect 831 876 835 880
rect 1079 879 1083 883
rect 1169 879 1173 883
rect 1040 875 1044 879
rect 1345 878 1349 882
rect 1435 878 1439 882
rect 1306 874 1310 878
rect -148 837 -144 841
rect -58 837 -54 841
rect 118 836 122 840
rect 208 836 212 840
rect 313 837 317 841
rect 529 843 533 847
rect 718 842 722 846
rect 1017 859 1021 863
rect 1099 858 1103 862
rect 1189 858 1193 862
rect 1283 858 1287 862
rect 1365 857 1369 861
rect 1455 857 1459 861
rect 834 847 838 851
rect 940 847 944 851
rect 394 830 398 834
rect -128 816 -124 820
rect 794 824 798 828
rect 854 826 858 830
rect 917 831 921 835
rect 1020 830 1024 834
rect 1286 829 1290 833
rect -38 816 -34 820
rect 138 815 142 819
rect 228 815 232 819
rect 371 814 375 818
rect 521 814 525 818
rect 1040 809 1044 813
rect 1306 808 1310 812
rect 920 802 924 806
rect 854 797 858 801
rect -189 776 -185 780
rect 374 785 378 789
rect 480 785 484 789
rect 831 781 835 785
rect 940 781 944 785
rect 1095 782 1099 786
rect 1185 782 1189 786
rect 1361 781 1365 785
rect 1451 781 1455 785
rect 334 762 338 766
rect 394 764 398 768
rect 457 769 461 773
rect 1072 766 1076 770
rect 1162 766 1166 770
rect -124 752 -120 756
rect -34 752 -30 756
rect 142 751 146 755
rect 232 751 236 755
rect 1338 765 1342 769
rect 1428 765 1432 769
rect 834 752 838 756
rect 460 740 464 744
rect -147 736 -143 740
rect -57 736 -53 740
rect 119 735 123 739
rect 209 735 213 739
rect 394 735 398 739
rect 854 731 858 735
rect 1075 737 1079 741
rect 1165 737 1169 741
rect 1341 736 1345 740
rect 1431 736 1435 740
rect 371 719 375 723
rect 480 719 484 723
rect -144 707 -140 711
rect -54 707 -50 711
rect 1095 716 1099 720
rect 1185 716 1189 720
rect 1361 715 1365 719
rect 1451 715 1455 719
rect -183 703 -179 707
rect 122 706 126 710
rect 212 706 216 710
rect 83 702 87 706
rect -206 687 -202 691
rect -124 686 -120 690
rect -34 686 -30 690
rect 60 686 64 690
rect 142 685 146 689
rect 232 685 236 689
rect 374 690 378 694
rect -203 658 -199 662
rect 394 669 398 673
rect 773 666 777 670
rect 1034 676 1038 680
rect 63 657 67 661
rect 854 659 858 663
rect 1099 652 1103 656
rect 1189 652 1193 656
rect 1365 651 1369 655
rect -183 637 -179 641
rect 831 643 835 647
rect 1455 651 1459 655
rect 83 636 87 640
rect 1076 636 1080 640
rect 1166 636 1170 640
rect 1342 635 1346 639
rect 1432 635 1436 639
rect 349 622 353 626
rect -128 610 -124 614
rect -38 610 -34 614
rect 138 609 142 613
rect 228 609 232 613
rect 834 614 838 618
rect 940 614 944 618
rect 326 606 330 610
rect 1079 607 1083 611
rect 1169 607 1173 611
rect 1040 603 1044 607
rect 1345 606 1349 610
rect 1435 606 1439 610
rect -151 594 -147 598
rect -61 594 -57 598
rect 115 593 119 597
rect 205 593 209 597
rect 390 591 394 595
rect 794 591 798 595
rect 854 593 858 597
rect 917 598 921 602
rect 1306 602 1310 606
rect 1017 587 1021 591
rect 329 577 333 581
rect -148 565 -144 569
rect -58 565 -54 569
rect 1099 586 1103 590
rect 1189 586 1193 590
rect 1283 586 1287 590
rect 1365 585 1369 589
rect 1455 585 1459 589
rect 118 564 122 568
rect 208 564 212 568
rect 920 569 924 573
rect 854 564 858 568
rect 349 556 353 560
rect 1020 558 1024 562
rect 1286 557 1290 561
rect -128 544 -124 548
rect -38 544 -34 548
rect 138 543 142 547
rect 228 543 232 547
rect 831 548 835 552
rect 940 548 944 552
rect 1040 537 1044 541
rect 1306 536 1310 540
rect -189 504 -185 508
rect 834 519 838 523
rect 313 502 317 506
rect 1095 510 1099 514
rect 1185 510 1189 514
rect 1361 509 1365 513
rect 394 495 398 499
rect 854 498 858 502
rect 1451 509 1455 513
rect 1072 494 1076 498
rect 1162 494 1166 498
rect 1338 493 1342 497
rect 1428 493 1432 497
rect -124 480 -120 484
rect -34 480 -30 484
rect 142 479 146 483
rect 232 479 236 483
rect 371 479 375 483
rect -147 464 -143 468
rect -57 464 -53 468
rect 119 463 123 467
rect 209 463 213 467
rect 1075 465 1079 469
rect 1165 465 1169 469
rect 1341 464 1345 468
rect 1431 464 1435 468
rect 374 450 378 454
rect 480 450 484 454
rect -144 435 -140 439
rect -54 435 -50 439
rect 1095 444 1099 448
rect 1185 444 1189 448
rect 1361 443 1365 447
rect 1451 443 1455 447
rect -183 431 -179 435
rect 122 434 126 438
rect 212 434 216 438
rect 83 430 87 434
rect 334 427 338 431
rect 394 429 398 433
rect 457 434 461 438
rect -206 415 -202 419
rect -124 414 -120 418
rect -34 414 -30 418
rect 60 414 64 418
rect 142 413 146 417
rect 232 413 236 417
rect 460 405 464 409
rect 1034 404 1038 408
rect 394 400 398 404
rect -203 386 -199 390
rect 63 385 67 389
rect 371 384 375 388
rect 480 384 484 388
rect 1099 380 1103 384
rect 1189 380 1193 384
rect 1365 379 1369 383
rect -183 365 -179 369
rect 1455 379 1459 383
rect 83 364 87 368
rect 1076 364 1080 368
rect 1166 364 1170 368
rect 374 355 378 359
rect 1342 363 1346 367
rect 1432 363 1436 367
rect -128 338 -124 342
rect -38 338 -34 342
rect 138 337 142 341
rect 228 337 232 341
rect 394 334 398 338
rect 1079 335 1083 339
rect 1169 335 1173 339
rect 1040 331 1044 335
rect 1345 334 1349 338
rect 1435 334 1439 338
rect 1306 330 1310 334
rect -151 322 -147 326
rect -61 322 -57 326
rect 115 321 119 325
rect 205 321 209 325
rect 1017 315 1021 319
rect 1099 314 1103 318
rect 1189 314 1193 318
rect 1283 314 1287 318
rect 1365 313 1369 317
rect 1455 313 1459 317
rect -148 293 -144 297
rect -58 293 -54 297
rect 118 292 122 296
rect 208 292 212 296
rect 349 287 353 291
rect 1020 286 1024 290
rect 1286 285 1290 289
rect -128 272 -124 276
rect -38 272 -34 276
rect 138 271 142 275
rect 228 271 232 275
rect 326 271 330 275
rect 390 256 394 260
rect 1040 265 1044 269
rect 1306 264 1310 268
rect -189 232 -185 236
rect 329 242 333 246
rect 349 221 353 225
rect -124 208 -120 212
rect -34 208 -30 212
rect 142 207 146 211
rect 232 207 236 211
rect -147 192 -143 196
rect -57 192 -53 196
rect 119 191 123 195
rect 209 191 213 195
rect -144 163 -140 167
rect -54 163 -50 167
rect -183 159 -179 163
rect 122 162 126 166
rect 212 162 216 166
rect 83 158 87 162
rect -206 143 -202 147
rect -124 142 -120 146
rect -34 142 -30 146
rect 60 142 64 146
rect 142 141 146 145
rect 232 141 236 145
rect -203 114 -199 118
rect 63 113 67 117
rect -183 93 -179 97
rect 83 92 87 96
rect -128 66 -124 70
rect -38 66 -34 70
rect 138 65 142 69
rect 228 65 232 69
rect -151 50 -147 54
rect -61 50 -57 54
rect 115 49 119 53
rect 205 49 209 53
rect -148 21 -144 25
rect -58 21 -54 25
rect 118 20 122 24
rect 208 20 212 24
rect -128 0 -124 4
rect -38 0 -34 4
rect 138 -1 142 3
rect 228 -1 232 3
rect -189 -40 -185 -36
rect -124 -64 -120 -60
rect -34 -64 -30 -60
rect 142 -65 146 -61
rect 232 -65 236 -61
rect -147 -80 -143 -76
rect -57 -80 -53 -76
rect 119 -81 123 -77
rect 209 -81 213 -77
rect -144 -109 -140 -105
rect -54 -109 -50 -105
rect -183 -113 -179 -109
rect 122 -110 126 -106
rect 212 -110 216 -106
rect 83 -114 87 -110
rect -206 -129 -202 -125
rect -124 -130 -120 -126
rect -34 -130 -30 -126
rect 60 -130 64 -126
rect 142 -131 146 -127
rect 232 -131 236 -127
rect -203 -158 -199 -154
rect 63 -159 67 -155
rect -183 -179 -179 -175
rect 83 -180 87 -176
<< metal1 >>
rect -236 1977 -124 1981
rect -92 1977 -34 1981
rect -236 1802 -232 1977
rect -151 1958 -147 1977
rect -128 1974 -124 1977
rect -104 1971 -100 1977
rect -109 1967 -100 1971
rect -173 1953 -169 1957
rect -173 1949 -163 1953
rect -173 1937 -169 1949
rect -155 1941 -141 1945
rect -117 1943 -109 1959
rect -104 1952 -100 1967
rect -92 1943 -88 1977
rect -61 1958 -57 1977
rect -38 1974 -34 1977
rect -14 1971 -10 1977
rect -19 1967 -10 1971
rect -117 1939 -88 1943
rect -83 1953 -79 1957
rect -83 1949 -73 1953
rect -117 1937 -109 1939
rect -83 1937 -79 1949
rect -65 1941 -51 1945
rect -27 1943 -19 1959
rect -14 1952 -10 1967
rect 30 1976 142 1980
rect 174 1976 232 1980
rect 30 1943 34 1976
rect 115 1957 119 1976
rect 138 1973 142 1976
rect 162 1970 166 1976
rect 157 1966 166 1970
rect -27 1939 34 1943
rect -27 1937 -19 1939
rect -133 1933 -109 1937
rect -43 1933 -19 1937
rect -148 1900 -144 1925
rect -117 1919 -109 1933
rect -104 1911 -100 1926
rect -109 1907 -100 1911
rect -128 1900 -124 1904
rect -104 1901 -100 1907
rect -148 1896 -124 1900
rect -58 1900 -54 1925
rect -27 1919 -19 1933
rect -14 1911 -10 1926
rect -19 1907 -10 1911
rect -38 1900 -34 1904
rect -14 1901 -10 1907
rect -58 1896 -34 1900
rect -188 1888 -164 1892
rect -182 1883 -178 1888
rect -174 1868 -170 1875
rect -148 1868 -144 1896
rect -58 1887 -54 1896
rect -58 1883 6 1887
rect -193 1864 -189 1868
rect -174 1864 -143 1868
rect -174 1863 -170 1864
rect -182 1850 -178 1855
rect -147 1851 -143 1864
rect -186 1846 -166 1850
rect -147 1847 -120 1851
rect -88 1848 -30 1851
rect -147 1828 -143 1847
rect -124 1844 -120 1847
rect -100 1841 -96 1847
rect -105 1837 -96 1841
rect -169 1823 -165 1827
rect -169 1819 -159 1823
rect -169 1807 -165 1819
rect -151 1811 -137 1815
rect -113 1813 -105 1829
rect -100 1822 -96 1837
rect -88 1813 -84 1848
rect -57 1847 -30 1848
rect -57 1828 -53 1847
rect -34 1844 -30 1847
rect -10 1841 -6 1847
rect -15 1837 -6 1841
rect -113 1809 -84 1813
rect -79 1823 -75 1827
rect -79 1819 -69 1823
rect -113 1807 -105 1809
rect -79 1807 -75 1819
rect -61 1811 -47 1815
rect -23 1813 -15 1829
rect -10 1822 -6 1837
rect 2 1813 6 1883
rect -23 1809 6 1813
rect -23 1807 -15 1809
rect -129 1803 -105 1807
rect -39 1803 -15 1807
rect -236 1798 -179 1802
rect -236 1721 -232 1798
rect -206 1779 -202 1798
rect -183 1795 -179 1798
rect -159 1792 -155 1798
rect -164 1788 -155 1792
rect -228 1774 -224 1778
rect -228 1770 -218 1774
rect -228 1758 -224 1770
rect -210 1762 -196 1766
rect -172 1764 -164 1780
rect -159 1773 -155 1788
rect -144 1770 -140 1795
rect -113 1789 -105 1803
rect -100 1781 -96 1796
rect -105 1777 -96 1781
rect -124 1770 -120 1774
rect -100 1771 -96 1777
rect -144 1766 -120 1770
rect -54 1770 -50 1795
rect -23 1789 -15 1803
rect -10 1781 -6 1796
rect -15 1777 -6 1781
rect -34 1770 -30 1774
rect -10 1771 -6 1777
rect -54 1766 -30 1770
rect -144 1764 -140 1766
rect -172 1760 -140 1764
rect -172 1758 -164 1760
rect -188 1754 -164 1758
rect -203 1721 -199 1746
rect -172 1740 -164 1754
rect -54 1757 -50 1766
rect 18 1757 22 1939
rect -54 1753 22 1757
rect 30 1801 34 1939
rect 93 1952 97 1956
rect 93 1948 103 1952
rect 93 1936 97 1948
rect 111 1940 125 1944
rect 149 1942 157 1958
rect 162 1951 166 1966
rect 174 1942 178 1976
rect 205 1957 209 1976
rect 228 1973 232 1976
rect 252 1970 256 1976
rect 247 1966 256 1970
rect 149 1938 178 1942
rect 183 1952 187 1956
rect 183 1948 193 1952
rect 149 1936 157 1938
rect 183 1936 187 1948
rect 201 1940 215 1944
rect 239 1942 247 1958
rect 252 1951 256 1966
rect 239 1938 288 1942
rect 239 1936 247 1938
rect 133 1932 157 1936
rect 223 1932 247 1936
rect 118 1899 122 1924
rect 149 1918 157 1932
rect 162 1910 166 1925
rect 157 1906 166 1910
rect 138 1899 142 1903
rect 162 1900 166 1906
rect 118 1895 142 1899
rect 208 1899 212 1924
rect 239 1918 247 1932
rect 252 1910 256 1925
rect 247 1906 256 1910
rect 228 1899 232 1903
rect 252 1900 256 1906
rect 208 1895 232 1899
rect 118 1867 122 1895
rect 208 1886 212 1895
rect 208 1882 272 1886
rect 114 1863 123 1867
rect 119 1850 123 1863
rect 119 1846 146 1850
rect 178 1847 236 1850
rect 119 1827 123 1846
rect 142 1843 146 1846
rect 166 1840 170 1846
rect 161 1836 170 1840
rect 97 1822 101 1826
rect 97 1818 107 1822
rect 97 1806 101 1818
rect 115 1810 129 1814
rect 153 1812 161 1828
rect 166 1821 170 1836
rect 178 1812 182 1847
rect 209 1846 236 1847
rect 209 1827 213 1846
rect 232 1843 236 1846
rect 256 1840 260 1846
rect 251 1836 260 1840
rect 153 1808 182 1812
rect 187 1822 191 1826
rect 187 1818 197 1822
rect 153 1806 161 1808
rect 187 1806 191 1818
rect 205 1810 219 1814
rect 243 1812 251 1828
rect 256 1821 260 1836
rect 268 1812 272 1882
rect 243 1808 272 1812
rect 243 1806 251 1808
rect 137 1802 161 1806
rect 227 1802 251 1806
rect 30 1797 87 1801
rect -159 1732 -155 1747
rect -164 1728 -155 1732
rect -183 1721 -179 1725
rect -159 1722 -155 1728
rect -236 1717 -179 1721
rect 30 1720 34 1797
rect 60 1778 64 1797
rect 83 1794 87 1797
rect 107 1791 111 1797
rect 102 1787 111 1791
rect 38 1773 42 1777
rect 38 1769 48 1773
rect 38 1757 42 1769
rect 56 1761 70 1765
rect 94 1763 102 1779
rect 107 1772 111 1787
rect 122 1769 126 1794
rect 153 1788 161 1802
rect 166 1780 170 1795
rect 161 1776 170 1780
rect 142 1769 146 1773
rect 166 1770 170 1776
rect 122 1765 146 1769
rect 212 1769 216 1794
rect 243 1788 251 1802
rect 256 1780 260 1795
rect 251 1776 260 1780
rect 232 1769 236 1773
rect 256 1770 260 1776
rect 212 1765 236 1769
rect 122 1763 126 1765
rect 94 1759 126 1763
rect 94 1757 102 1759
rect 78 1753 102 1757
rect 63 1720 67 1745
rect 94 1739 102 1753
rect 212 1756 216 1765
rect 284 1756 288 1938
rect 212 1752 288 1756
rect 107 1731 111 1746
rect 102 1727 111 1731
rect 83 1720 87 1724
rect 107 1721 111 1727
rect 30 1716 87 1720
rect -236 1705 -124 1709
rect -92 1705 -34 1709
rect -236 1530 -232 1705
rect -151 1686 -147 1705
rect -128 1702 -124 1705
rect -104 1699 -100 1705
rect -109 1695 -100 1699
rect -173 1681 -169 1685
rect -173 1677 -163 1681
rect -173 1665 -169 1677
rect -155 1669 -141 1673
rect -117 1671 -109 1687
rect -104 1680 -100 1695
rect -92 1671 -88 1705
rect -61 1686 -57 1705
rect -38 1702 -34 1705
rect -14 1699 -10 1705
rect -19 1695 -10 1699
rect -117 1667 -88 1671
rect -83 1681 -79 1685
rect -83 1677 -73 1681
rect -117 1665 -109 1667
rect -83 1665 -79 1677
rect -65 1669 -51 1673
rect -27 1671 -19 1687
rect -14 1680 -10 1695
rect 30 1704 142 1708
rect 174 1704 232 1708
rect 30 1671 34 1704
rect 115 1685 119 1704
rect 138 1701 142 1704
rect 162 1698 166 1704
rect 157 1694 166 1698
rect -27 1667 34 1671
rect -27 1665 -19 1667
rect -133 1661 -109 1665
rect -43 1661 -19 1665
rect -148 1628 -144 1653
rect -117 1647 -109 1661
rect -104 1639 -100 1654
rect -109 1635 -100 1639
rect -128 1628 -124 1632
rect -104 1629 -100 1635
rect -148 1624 -124 1628
rect -58 1628 -54 1653
rect -27 1647 -19 1661
rect -14 1639 -10 1654
rect -19 1635 -10 1639
rect -38 1628 -34 1632
rect -14 1629 -10 1635
rect -58 1624 -34 1628
rect -188 1616 -164 1620
rect -182 1611 -178 1616
rect -174 1596 -170 1603
rect -148 1596 -144 1624
rect -58 1615 -54 1624
rect -58 1611 6 1615
rect -193 1592 -189 1596
rect -174 1592 -143 1596
rect -174 1591 -170 1592
rect -182 1578 -178 1583
rect -147 1579 -143 1592
rect -186 1574 -166 1578
rect -147 1575 -120 1579
rect -88 1576 -30 1579
rect -147 1556 -143 1575
rect -124 1572 -120 1575
rect -100 1569 -96 1575
rect -105 1565 -96 1569
rect -169 1551 -165 1555
rect -169 1547 -159 1551
rect -169 1535 -165 1547
rect -151 1539 -137 1543
rect -113 1541 -105 1557
rect -100 1550 -96 1565
rect -88 1541 -84 1576
rect -57 1575 -30 1576
rect -57 1556 -53 1575
rect -34 1572 -30 1575
rect -10 1569 -6 1575
rect -15 1565 -6 1569
rect -113 1537 -84 1541
rect -79 1551 -75 1555
rect -79 1547 -69 1551
rect -113 1535 -105 1537
rect -79 1535 -75 1547
rect -61 1539 -47 1543
rect -23 1541 -15 1557
rect -10 1550 -6 1565
rect 2 1541 6 1611
rect -23 1537 6 1541
rect -23 1535 -15 1537
rect -129 1531 -105 1535
rect -39 1531 -15 1535
rect -236 1526 -179 1530
rect -236 1449 -232 1526
rect -206 1507 -202 1526
rect -183 1523 -179 1526
rect -159 1520 -155 1526
rect -164 1516 -155 1520
rect -228 1502 -224 1506
rect -228 1498 -218 1502
rect -228 1486 -224 1498
rect -210 1490 -196 1494
rect -172 1492 -164 1508
rect -159 1501 -155 1516
rect -144 1498 -140 1523
rect -113 1517 -105 1531
rect -100 1509 -96 1524
rect -105 1505 -96 1509
rect -124 1498 -120 1502
rect -100 1499 -96 1505
rect -144 1494 -120 1498
rect -54 1498 -50 1523
rect -23 1517 -15 1531
rect -10 1509 -6 1524
rect -15 1505 -6 1509
rect -34 1498 -30 1502
rect -10 1499 -6 1505
rect -54 1494 -30 1498
rect -144 1492 -140 1494
rect -172 1488 -140 1492
rect -172 1486 -164 1488
rect -188 1482 -164 1486
rect -203 1449 -199 1474
rect -172 1468 -164 1482
rect -54 1485 -50 1494
rect 18 1485 22 1667
rect -54 1481 22 1485
rect 30 1529 34 1667
rect 93 1680 97 1684
rect 93 1676 103 1680
rect 93 1664 97 1676
rect 111 1668 125 1672
rect 149 1670 157 1686
rect 162 1679 166 1694
rect 174 1670 178 1704
rect 205 1685 209 1704
rect 228 1701 232 1704
rect 252 1698 256 1704
rect 247 1694 256 1698
rect 149 1666 178 1670
rect 183 1680 187 1684
rect 183 1676 193 1680
rect 149 1664 157 1666
rect 183 1664 187 1676
rect 201 1668 215 1672
rect 239 1670 247 1686
rect 252 1679 256 1694
rect 239 1666 288 1670
rect 239 1664 247 1666
rect 133 1660 157 1664
rect 223 1660 247 1664
rect 118 1627 122 1652
rect 149 1646 157 1660
rect 162 1638 166 1653
rect 157 1634 166 1638
rect 138 1627 142 1631
rect 162 1628 166 1634
rect 118 1623 142 1627
rect 208 1627 212 1652
rect 239 1646 247 1660
rect 252 1638 256 1653
rect 247 1634 256 1638
rect 228 1627 232 1631
rect 252 1628 256 1634
rect 208 1623 232 1627
rect 118 1595 122 1623
rect 208 1614 212 1623
rect 208 1610 272 1614
rect 114 1591 123 1595
rect 119 1578 123 1591
rect 119 1574 146 1578
rect 178 1575 236 1578
rect 119 1555 123 1574
rect 142 1571 146 1574
rect 166 1568 170 1574
rect 161 1564 170 1568
rect 97 1550 101 1554
rect 97 1546 107 1550
rect 97 1534 101 1546
rect 115 1538 129 1542
rect 153 1540 161 1556
rect 166 1549 170 1564
rect 178 1540 182 1575
rect 209 1574 236 1575
rect 209 1555 213 1574
rect 232 1571 236 1574
rect 256 1568 260 1574
rect 251 1564 260 1568
rect 153 1536 182 1540
rect 187 1550 191 1554
rect 187 1546 197 1550
rect 153 1534 161 1536
rect 187 1534 191 1546
rect 205 1538 219 1542
rect 243 1540 251 1556
rect 256 1549 260 1564
rect 268 1540 272 1610
rect 243 1536 272 1540
rect 243 1534 251 1536
rect 137 1530 161 1534
rect 227 1530 251 1534
rect 30 1525 87 1529
rect -159 1460 -155 1475
rect -164 1456 -155 1460
rect -183 1449 -179 1453
rect -159 1450 -155 1456
rect -236 1445 -179 1449
rect 30 1448 34 1525
rect 60 1506 64 1525
rect 83 1522 87 1525
rect 107 1519 111 1525
rect 102 1515 111 1519
rect 38 1501 42 1505
rect 38 1497 48 1501
rect 38 1485 42 1497
rect 56 1489 70 1493
rect 94 1491 102 1507
rect 107 1500 111 1515
rect 122 1497 126 1522
rect 153 1516 161 1530
rect 166 1508 170 1523
rect 161 1504 170 1508
rect 142 1497 146 1501
rect 166 1498 170 1504
rect 122 1493 146 1497
rect 212 1497 216 1522
rect 243 1516 251 1530
rect 256 1508 260 1523
rect 251 1504 260 1508
rect 232 1497 236 1501
rect 256 1498 260 1504
rect 212 1493 236 1497
rect 122 1491 126 1493
rect 94 1487 126 1491
rect 94 1485 102 1487
rect 78 1481 102 1485
rect 63 1448 67 1473
rect 94 1467 102 1481
rect 212 1484 216 1493
rect 284 1484 288 1666
rect 987 1605 1099 1609
rect 1131 1605 1189 1609
rect 314 1531 338 1535
rect 320 1526 324 1531
rect 328 1511 332 1518
rect 212 1480 288 1484
rect 304 1507 313 1511
rect 328 1507 398 1511
rect 107 1459 111 1474
rect 102 1455 111 1459
rect 83 1448 87 1452
rect 107 1449 111 1455
rect 30 1444 87 1448
rect -236 1433 -124 1437
rect -92 1433 -34 1437
rect -236 1258 -232 1433
rect -151 1414 -147 1433
rect -128 1430 -124 1433
rect -104 1427 -100 1433
rect -109 1423 -100 1427
rect -173 1409 -169 1413
rect -173 1405 -163 1409
rect -173 1393 -169 1405
rect -155 1397 -141 1401
rect -117 1399 -109 1415
rect -104 1408 -100 1423
rect -92 1399 -88 1433
rect -61 1414 -57 1433
rect -38 1430 -34 1433
rect -14 1427 -10 1433
rect -19 1423 -10 1427
rect -117 1395 -88 1399
rect -83 1409 -79 1413
rect -83 1405 -73 1409
rect -117 1393 -109 1395
rect -83 1393 -79 1405
rect -65 1397 -51 1401
rect -27 1399 -19 1415
rect -14 1408 -10 1423
rect 30 1432 142 1436
rect 174 1432 232 1436
rect 30 1399 34 1432
rect 115 1413 119 1432
rect 138 1429 142 1432
rect 162 1426 166 1432
rect 157 1422 166 1426
rect -27 1395 34 1399
rect -27 1393 -19 1395
rect -133 1389 -109 1393
rect -43 1389 -19 1393
rect -148 1356 -144 1381
rect -117 1375 -109 1389
rect -104 1367 -100 1382
rect -109 1363 -100 1367
rect -128 1356 -124 1360
rect -104 1357 -100 1363
rect -148 1352 -124 1356
rect -58 1356 -54 1381
rect -27 1375 -19 1389
rect -14 1367 -10 1382
rect -19 1363 -10 1367
rect -38 1356 -34 1360
rect -14 1357 -10 1363
rect -58 1352 -34 1356
rect -188 1344 -164 1348
rect -182 1339 -178 1344
rect -174 1324 -170 1331
rect -148 1324 -144 1352
rect -58 1343 -54 1352
rect -58 1339 6 1343
rect -193 1320 -189 1324
rect -174 1320 -143 1324
rect -174 1319 -170 1320
rect -182 1306 -178 1311
rect -147 1307 -143 1320
rect -186 1302 -166 1306
rect -147 1303 -120 1307
rect -88 1304 -30 1307
rect -147 1284 -143 1303
rect -124 1300 -120 1303
rect -100 1297 -96 1303
rect -105 1293 -96 1297
rect -169 1279 -165 1283
rect -169 1275 -159 1279
rect -169 1263 -165 1275
rect -151 1267 -137 1271
rect -113 1269 -105 1285
rect -100 1278 -96 1293
rect -88 1269 -84 1304
rect -57 1303 -30 1304
rect -57 1284 -53 1303
rect -34 1300 -30 1303
rect -10 1297 -6 1303
rect -15 1293 -6 1297
rect -113 1265 -84 1269
rect -79 1279 -75 1283
rect -79 1275 -69 1279
rect -113 1263 -105 1265
rect -79 1263 -75 1275
rect -61 1267 -47 1271
rect -23 1269 -15 1285
rect -10 1278 -6 1293
rect 2 1269 6 1339
rect -23 1265 6 1269
rect -23 1263 -15 1265
rect -129 1259 -105 1263
rect -39 1259 -15 1263
rect -236 1254 -179 1258
rect -236 1177 -232 1254
rect -206 1235 -202 1254
rect -183 1251 -179 1254
rect -159 1248 -155 1254
rect -164 1244 -155 1248
rect -228 1230 -224 1234
rect -228 1226 -218 1230
rect -228 1214 -224 1226
rect -210 1218 -196 1222
rect -172 1220 -164 1236
rect -159 1229 -155 1244
rect -144 1226 -140 1251
rect -113 1245 -105 1259
rect -100 1237 -96 1252
rect -105 1233 -96 1237
rect -124 1226 -120 1230
rect -100 1227 -96 1233
rect -144 1222 -120 1226
rect -54 1226 -50 1251
rect -23 1245 -15 1259
rect -10 1237 -6 1252
rect -15 1233 -6 1237
rect -34 1226 -30 1230
rect -10 1227 -6 1233
rect -54 1222 -30 1226
rect -144 1220 -140 1222
rect -172 1216 -140 1220
rect -172 1214 -164 1216
rect -188 1210 -164 1214
rect -203 1177 -199 1202
rect -172 1196 -164 1210
rect -54 1213 -50 1222
rect 18 1213 22 1395
rect -54 1209 22 1213
rect 30 1257 34 1395
rect 93 1408 97 1412
rect 93 1404 103 1408
rect 93 1392 97 1404
rect 111 1396 125 1400
rect 149 1398 157 1414
rect 162 1407 166 1422
rect 174 1398 178 1432
rect 205 1413 209 1432
rect 228 1429 232 1432
rect 252 1426 256 1432
rect 247 1422 256 1426
rect 149 1394 178 1398
rect 183 1408 187 1412
rect 183 1404 193 1408
rect 149 1392 157 1394
rect 183 1392 187 1404
rect 201 1396 215 1400
rect 239 1398 247 1414
rect 252 1407 256 1422
rect 239 1394 288 1398
rect 239 1392 247 1394
rect 133 1388 157 1392
rect 223 1388 247 1392
rect 118 1355 122 1380
rect 149 1374 157 1388
rect 162 1366 166 1381
rect 157 1362 166 1366
rect 138 1355 142 1359
rect 162 1356 166 1362
rect 118 1351 142 1355
rect 208 1355 212 1380
rect 239 1374 247 1388
rect 252 1366 256 1381
rect 247 1362 256 1366
rect 228 1355 232 1359
rect 252 1356 256 1362
rect 208 1351 232 1355
rect 118 1323 122 1351
rect 208 1342 212 1351
rect 208 1338 272 1342
rect 114 1319 123 1323
rect 119 1306 123 1319
rect 119 1302 146 1306
rect 178 1303 236 1306
rect 119 1283 123 1302
rect 142 1299 146 1302
rect 166 1296 170 1302
rect 161 1292 170 1296
rect 97 1278 101 1282
rect 97 1274 107 1278
rect 97 1262 101 1274
rect 115 1266 129 1270
rect 153 1268 161 1284
rect 166 1277 170 1292
rect 178 1268 182 1303
rect 209 1302 236 1303
rect 209 1283 213 1302
rect 232 1299 236 1302
rect 256 1296 260 1302
rect 251 1292 260 1296
rect 153 1264 182 1268
rect 187 1278 191 1282
rect 187 1274 197 1278
rect 153 1262 161 1264
rect 187 1262 191 1274
rect 205 1266 219 1270
rect 243 1268 251 1284
rect 256 1277 260 1292
rect 268 1268 272 1338
rect 243 1264 272 1268
rect 243 1262 251 1264
rect 137 1258 161 1262
rect 227 1258 251 1262
rect 30 1253 87 1257
rect -159 1188 -155 1203
rect -164 1184 -155 1188
rect -183 1177 -179 1181
rect -159 1178 -155 1184
rect -236 1173 -179 1177
rect 30 1176 34 1253
rect 60 1234 64 1253
rect 83 1250 87 1253
rect 107 1247 111 1253
rect 102 1243 111 1247
rect 38 1229 42 1233
rect 38 1225 48 1229
rect 38 1213 42 1225
rect 56 1217 70 1221
rect 94 1219 102 1235
rect 107 1228 111 1243
rect 122 1225 126 1250
rect 153 1244 161 1258
rect 166 1236 170 1251
rect 161 1232 170 1236
rect 142 1225 146 1229
rect 166 1226 170 1232
rect 122 1221 146 1225
rect 212 1225 216 1250
rect 243 1244 251 1258
rect 256 1236 260 1251
rect 251 1232 260 1236
rect 232 1225 236 1229
rect 256 1226 260 1232
rect 212 1221 236 1225
rect 122 1219 126 1221
rect 94 1215 126 1219
rect 94 1213 102 1215
rect 78 1209 102 1213
rect 63 1176 67 1201
rect 94 1195 102 1209
rect 212 1212 216 1221
rect 284 1212 288 1394
rect 304 1335 308 1507
rect 328 1506 332 1507
rect 320 1493 324 1498
rect 316 1489 336 1493
rect 371 1488 375 1507
rect 394 1504 398 1507
rect 418 1501 422 1507
rect 413 1497 422 1501
rect 349 1483 353 1487
rect 349 1479 359 1483
rect 349 1467 353 1479
rect 367 1471 381 1475
rect 405 1473 413 1489
rect 418 1482 422 1497
rect 405 1469 461 1473
rect 405 1467 413 1469
rect 389 1463 413 1467
rect 374 1444 378 1455
rect 405 1449 413 1463
rect 457 1466 461 1469
rect 457 1462 484 1466
rect 334 1440 378 1444
rect 418 1441 422 1456
rect 457 1443 461 1462
rect 480 1459 484 1462
rect 504 1456 508 1462
rect 499 1452 508 1456
rect 334 1436 338 1440
rect 316 1429 320 1433
rect 358 1429 362 1435
rect 316 1425 325 1429
rect 353 1425 362 1429
rect 374 1430 378 1440
rect 413 1437 422 1441
rect 394 1430 398 1434
rect 418 1431 422 1437
rect 435 1438 439 1442
rect 435 1434 445 1438
rect 374 1426 398 1430
rect 316 1413 320 1425
rect 333 1417 345 1421
rect 334 1406 338 1417
rect 358 1411 362 1425
rect 435 1422 439 1434
rect 453 1426 467 1430
rect 491 1428 499 1444
rect 504 1437 508 1452
rect 987 1430 991 1605
rect 1072 1586 1076 1605
rect 1095 1602 1099 1605
rect 1119 1599 1123 1605
rect 1114 1595 1123 1599
rect 1050 1581 1054 1585
rect 1050 1577 1060 1581
rect 1050 1565 1054 1577
rect 1068 1569 1082 1573
rect 1106 1571 1114 1587
rect 1119 1580 1123 1595
rect 1131 1571 1135 1605
rect 1162 1586 1166 1605
rect 1185 1602 1189 1605
rect 1209 1599 1213 1605
rect 1204 1595 1213 1599
rect 1106 1567 1135 1571
rect 1140 1581 1144 1585
rect 1140 1577 1150 1581
rect 1106 1565 1114 1567
rect 1140 1565 1144 1577
rect 1158 1569 1172 1573
rect 1196 1571 1204 1587
rect 1209 1580 1213 1595
rect 1253 1604 1365 1608
rect 1397 1604 1455 1608
rect 1253 1571 1257 1604
rect 1338 1585 1342 1604
rect 1361 1601 1365 1604
rect 1385 1598 1389 1604
rect 1380 1594 1389 1598
rect 1196 1567 1257 1571
rect 1196 1565 1204 1567
rect 1090 1561 1114 1565
rect 1180 1561 1204 1565
rect 1075 1528 1079 1553
rect 1106 1547 1114 1561
rect 1119 1539 1123 1554
rect 1114 1535 1123 1539
rect 1095 1528 1099 1532
rect 1119 1529 1123 1535
rect 1075 1524 1099 1528
rect 1165 1528 1169 1553
rect 1196 1547 1204 1561
rect 1209 1539 1213 1554
rect 1204 1535 1213 1539
rect 1185 1528 1189 1532
rect 1209 1529 1213 1535
rect 1165 1524 1189 1528
rect 1035 1516 1059 1520
rect 1041 1511 1045 1516
rect 1049 1496 1053 1503
rect 1075 1496 1079 1524
rect 1165 1515 1169 1524
rect 1165 1511 1229 1515
rect 1030 1492 1034 1496
rect 1049 1492 1080 1496
rect 1049 1491 1053 1492
rect 1041 1478 1045 1483
rect 1076 1479 1080 1492
rect 1037 1474 1057 1478
rect 1076 1475 1103 1479
rect 1135 1476 1193 1479
rect 1076 1456 1080 1475
rect 1099 1472 1103 1475
rect 1123 1469 1127 1475
rect 1118 1465 1127 1469
rect 1054 1451 1058 1455
rect 1054 1447 1064 1451
rect 1054 1435 1058 1447
rect 1072 1439 1086 1443
rect 1110 1441 1118 1457
rect 1123 1450 1127 1465
rect 1135 1441 1139 1476
rect 1166 1475 1193 1476
rect 1166 1456 1170 1475
rect 1189 1472 1193 1475
rect 1213 1469 1217 1475
rect 1208 1465 1217 1469
rect 1110 1437 1139 1441
rect 1144 1451 1148 1455
rect 1144 1447 1154 1451
rect 1110 1435 1118 1437
rect 1144 1435 1148 1447
rect 1162 1439 1176 1443
rect 1200 1441 1208 1457
rect 1213 1450 1217 1465
rect 1225 1441 1229 1511
rect 1200 1437 1229 1441
rect 1200 1435 1208 1437
rect 1094 1431 1118 1435
rect 1184 1431 1208 1435
rect 491 1424 514 1428
rect 987 1426 1044 1430
rect 491 1422 499 1424
rect 475 1418 499 1422
rect 371 1412 398 1416
rect 371 1406 375 1412
rect 334 1402 375 1406
rect 394 1409 398 1412
rect 418 1406 422 1412
rect 413 1402 422 1406
rect 371 1393 375 1402
rect 349 1388 353 1392
rect 349 1384 359 1388
rect 349 1372 353 1384
rect 367 1376 381 1380
rect 405 1378 413 1394
rect 418 1387 422 1402
rect 460 1385 464 1410
rect 491 1404 499 1418
rect 504 1396 508 1411
rect 499 1392 508 1396
rect 480 1385 484 1389
rect 504 1386 508 1392
rect 774 1389 798 1393
rect 460 1381 484 1385
rect 780 1384 784 1389
rect 460 1378 464 1381
rect 405 1374 464 1378
rect 405 1372 413 1374
rect 389 1368 413 1372
rect 788 1369 792 1376
rect 374 1335 378 1360
rect 405 1354 413 1368
rect 764 1365 773 1369
rect 788 1365 858 1369
rect 418 1346 422 1361
rect 413 1342 422 1346
rect 394 1335 398 1339
rect 418 1336 422 1342
rect 304 1331 398 1335
rect 326 1299 353 1303
rect 326 1280 330 1299
rect 349 1296 353 1299
rect 373 1293 377 1299
rect 368 1289 377 1293
rect 304 1275 308 1279
rect 304 1271 314 1275
rect 304 1259 308 1271
rect 322 1263 336 1267
rect 360 1265 368 1281
rect 373 1274 377 1289
rect 391 1285 415 1289
rect 397 1280 401 1285
rect 405 1265 409 1272
rect 360 1261 390 1265
rect 405 1261 426 1265
rect 360 1259 368 1261
rect 405 1260 409 1261
rect 344 1255 368 1259
rect 329 1222 333 1247
rect 360 1241 368 1255
rect 373 1233 377 1248
rect 397 1247 401 1252
rect 393 1243 413 1247
rect 368 1229 377 1233
rect 349 1222 353 1226
rect 373 1223 377 1229
rect 329 1218 353 1222
rect 212 1208 288 1212
rect 107 1187 111 1202
rect 314 1196 338 1200
rect 102 1183 111 1187
rect 320 1191 324 1196
rect 764 1193 768 1365
rect 788 1364 792 1365
rect 780 1351 784 1356
rect 776 1347 796 1351
rect 831 1346 835 1365
rect 854 1362 858 1365
rect 878 1359 882 1365
rect 873 1355 882 1359
rect 809 1341 813 1345
rect 809 1337 819 1341
rect 809 1325 813 1337
rect 827 1329 841 1333
rect 865 1331 873 1347
rect 878 1340 882 1355
rect 987 1349 991 1426
rect 1017 1407 1021 1426
rect 1040 1423 1044 1426
rect 1064 1420 1068 1426
rect 1059 1416 1068 1420
rect 995 1402 999 1406
rect 995 1398 1005 1402
rect 995 1386 999 1398
rect 1013 1390 1027 1394
rect 1051 1392 1059 1408
rect 1064 1401 1068 1416
rect 1079 1398 1083 1423
rect 1110 1417 1118 1431
rect 1123 1409 1127 1424
rect 1118 1405 1127 1409
rect 1099 1398 1103 1402
rect 1123 1399 1127 1405
rect 1079 1394 1103 1398
rect 1169 1398 1173 1423
rect 1200 1417 1208 1431
rect 1213 1409 1217 1424
rect 1208 1405 1217 1409
rect 1189 1398 1193 1402
rect 1213 1399 1217 1405
rect 1169 1394 1193 1398
rect 1079 1392 1083 1394
rect 1051 1388 1083 1392
rect 1051 1386 1059 1388
rect 1035 1382 1059 1386
rect 1020 1349 1024 1374
rect 1051 1368 1059 1382
rect 1169 1385 1173 1394
rect 1241 1385 1245 1567
rect 1169 1381 1245 1385
rect 1253 1429 1257 1567
rect 1316 1580 1320 1584
rect 1316 1576 1326 1580
rect 1316 1564 1320 1576
rect 1334 1568 1348 1572
rect 1372 1570 1380 1586
rect 1385 1579 1389 1594
rect 1397 1570 1401 1604
rect 1428 1585 1432 1604
rect 1451 1601 1455 1604
rect 1475 1598 1479 1604
rect 1470 1594 1479 1598
rect 1372 1566 1401 1570
rect 1406 1580 1410 1584
rect 1406 1576 1416 1580
rect 1372 1564 1380 1566
rect 1406 1564 1410 1576
rect 1424 1568 1438 1572
rect 1462 1570 1470 1586
rect 1475 1579 1479 1594
rect 1462 1566 1511 1570
rect 1462 1564 1470 1566
rect 1356 1560 1380 1564
rect 1446 1560 1470 1564
rect 1341 1527 1345 1552
rect 1372 1546 1380 1560
rect 1385 1538 1389 1553
rect 1380 1534 1389 1538
rect 1361 1527 1365 1531
rect 1385 1528 1389 1534
rect 1341 1523 1365 1527
rect 1431 1527 1435 1552
rect 1462 1546 1470 1560
rect 1475 1538 1479 1553
rect 1470 1534 1479 1538
rect 1451 1527 1455 1531
rect 1475 1528 1479 1534
rect 1431 1523 1455 1527
rect 1341 1495 1345 1523
rect 1431 1514 1435 1523
rect 1431 1510 1495 1514
rect 1337 1491 1346 1495
rect 1342 1478 1346 1491
rect 1342 1474 1369 1478
rect 1401 1475 1459 1478
rect 1342 1455 1346 1474
rect 1365 1471 1369 1474
rect 1389 1468 1393 1474
rect 1384 1464 1393 1468
rect 1320 1450 1324 1454
rect 1320 1446 1330 1450
rect 1320 1434 1324 1446
rect 1338 1438 1352 1442
rect 1376 1440 1384 1456
rect 1389 1449 1393 1464
rect 1401 1440 1405 1475
rect 1432 1474 1459 1475
rect 1432 1455 1436 1474
rect 1455 1471 1459 1474
rect 1479 1468 1483 1474
rect 1474 1464 1483 1468
rect 1376 1436 1405 1440
rect 1410 1450 1414 1454
rect 1410 1446 1420 1450
rect 1376 1434 1384 1436
rect 1410 1434 1414 1446
rect 1428 1438 1442 1442
rect 1466 1440 1474 1456
rect 1479 1449 1483 1464
rect 1491 1440 1495 1510
rect 1466 1436 1495 1440
rect 1466 1434 1474 1436
rect 1360 1430 1384 1434
rect 1450 1430 1474 1434
rect 1253 1425 1310 1429
rect 1064 1360 1068 1375
rect 1059 1356 1068 1360
rect 1040 1349 1044 1353
rect 1064 1350 1068 1356
rect 987 1345 1044 1349
rect 1253 1348 1257 1425
rect 1283 1406 1287 1425
rect 1306 1422 1310 1425
rect 1330 1419 1334 1425
rect 1325 1415 1334 1419
rect 1261 1401 1265 1405
rect 1261 1397 1271 1401
rect 1261 1385 1265 1397
rect 1279 1389 1293 1393
rect 1317 1391 1325 1407
rect 1330 1400 1334 1415
rect 1345 1397 1349 1422
rect 1376 1416 1384 1430
rect 1389 1408 1393 1423
rect 1384 1404 1393 1408
rect 1365 1397 1369 1401
rect 1389 1398 1393 1404
rect 1345 1393 1369 1397
rect 1435 1397 1439 1422
rect 1466 1416 1474 1430
rect 1479 1408 1483 1423
rect 1474 1404 1483 1408
rect 1455 1397 1459 1401
rect 1479 1398 1483 1404
rect 1435 1393 1459 1397
rect 1345 1391 1349 1393
rect 1317 1387 1349 1391
rect 1317 1385 1325 1387
rect 1301 1381 1325 1385
rect 1286 1348 1290 1373
rect 1317 1367 1325 1381
rect 1435 1384 1439 1393
rect 1507 1384 1511 1566
rect 1435 1380 1511 1384
rect 1330 1359 1334 1374
rect 1325 1355 1334 1359
rect 1306 1348 1310 1352
rect 1330 1349 1334 1355
rect 1253 1344 1310 1348
rect 987 1333 1099 1337
rect 1131 1333 1189 1337
rect 865 1327 921 1331
rect 865 1325 873 1327
rect 849 1321 873 1325
rect 834 1302 838 1313
rect 865 1307 873 1321
rect 917 1324 921 1327
rect 917 1320 944 1324
rect 794 1298 838 1302
rect 878 1299 882 1314
rect 917 1301 921 1320
rect 940 1317 944 1320
rect 964 1314 968 1320
rect 959 1310 968 1314
rect 794 1294 798 1298
rect 776 1287 780 1291
rect 818 1287 822 1293
rect 776 1283 785 1287
rect 813 1283 822 1287
rect 834 1288 838 1298
rect 873 1295 882 1299
rect 854 1288 858 1292
rect 878 1289 882 1295
rect 895 1296 899 1300
rect 895 1292 905 1296
rect 834 1284 858 1288
rect 776 1271 780 1283
rect 793 1275 805 1279
rect 794 1264 798 1275
rect 818 1269 822 1283
rect 895 1280 899 1292
rect 913 1284 927 1288
rect 951 1286 959 1302
rect 964 1295 968 1310
rect 951 1282 971 1286
rect 951 1280 959 1282
rect 935 1276 959 1280
rect 831 1270 858 1274
rect 831 1264 835 1270
rect 794 1260 835 1264
rect 854 1267 858 1270
rect 878 1264 882 1270
rect 873 1260 882 1264
rect 831 1251 835 1260
rect 809 1246 813 1250
rect 809 1242 819 1246
rect 809 1230 813 1242
rect 827 1234 841 1238
rect 865 1236 873 1252
rect 878 1245 882 1260
rect 920 1243 924 1268
rect 951 1262 959 1276
rect 964 1254 968 1269
rect 959 1250 968 1254
rect 940 1243 944 1247
rect 964 1244 968 1250
rect 920 1239 944 1243
rect 920 1236 924 1239
rect 865 1232 924 1236
rect 865 1230 873 1232
rect 849 1226 873 1230
rect 834 1193 838 1218
rect 865 1212 873 1226
rect 878 1204 882 1219
rect 873 1200 882 1204
rect 854 1193 858 1197
rect 878 1194 882 1200
rect 764 1189 858 1193
rect 83 1176 87 1180
rect 107 1177 111 1183
rect 328 1176 332 1183
rect 30 1172 87 1176
rect 304 1172 313 1176
rect 328 1172 398 1176
rect -236 1161 -124 1165
rect -92 1161 -34 1165
rect -236 986 -232 1161
rect -151 1142 -147 1161
rect -128 1158 -124 1161
rect -104 1155 -100 1161
rect -109 1151 -100 1155
rect -173 1137 -169 1141
rect -173 1133 -163 1137
rect -173 1121 -169 1133
rect -155 1125 -141 1129
rect -117 1127 -109 1143
rect -104 1136 -100 1151
rect -92 1127 -88 1161
rect -61 1142 -57 1161
rect -38 1158 -34 1161
rect -14 1155 -10 1161
rect -19 1151 -10 1155
rect -117 1123 -88 1127
rect -83 1137 -79 1141
rect -83 1133 -73 1137
rect -117 1121 -109 1123
rect -83 1121 -79 1133
rect -65 1125 -51 1129
rect -27 1127 -19 1143
rect -14 1136 -10 1151
rect 30 1160 142 1164
rect 174 1160 232 1164
rect 30 1127 34 1160
rect 115 1141 119 1160
rect 138 1157 142 1160
rect 162 1154 166 1160
rect 157 1150 166 1154
rect -27 1123 34 1127
rect -27 1121 -19 1123
rect -133 1117 -109 1121
rect -43 1117 -19 1121
rect -148 1084 -144 1109
rect -117 1103 -109 1117
rect -104 1095 -100 1110
rect -109 1091 -100 1095
rect -128 1084 -124 1088
rect -104 1085 -100 1091
rect -148 1080 -124 1084
rect -58 1084 -54 1109
rect -27 1103 -19 1117
rect -14 1095 -10 1110
rect -19 1091 -10 1095
rect -38 1084 -34 1088
rect -14 1085 -10 1091
rect -58 1080 -34 1084
rect -188 1072 -164 1076
rect -182 1067 -178 1072
rect -174 1052 -170 1059
rect -148 1052 -144 1080
rect -58 1071 -54 1080
rect -58 1067 6 1071
rect -193 1048 -189 1052
rect -174 1048 -143 1052
rect -174 1047 -170 1048
rect -182 1034 -178 1039
rect -147 1035 -143 1048
rect -186 1030 -166 1034
rect -147 1031 -120 1035
rect -88 1032 -30 1035
rect -147 1012 -143 1031
rect -124 1028 -120 1031
rect -100 1025 -96 1031
rect -105 1021 -96 1025
rect -169 1007 -165 1011
rect -169 1003 -159 1007
rect -169 991 -165 1003
rect -151 995 -137 999
rect -113 997 -105 1013
rect -100 1006 -96 1021
rect -88 997 -84 1032
rect -57 1031 -30 1032
rect -57 1012 -53 1031
rect -34 1028 -30 1031
rect -10 1025 -6 1031
rect -15 1021 -6 1025
rect -113 993 -84 997
rect -79 1007 -75 1011
rect -79 1003 -69 1007
rect -113 991 -105 993
rect -79 991 -75 1003
rect -61 995 -47 999
rect -23 997 -15 1013
rect -10 1006 -6 1021
rect 2 997 6 1067
rect -23 993 6 997
rect -23 991 -15 993
rect -129 987 -105 991
rect -39 987 -15 991
rect -236 982 -179 986
rect -236 905 -232 982
rect -206 963 -202 982
rect -183 979 -179 982
rect -159 976 -155 982
rect -164 972 -155 976
rect -228 958 -224 962
rect -228 954 -218 958
rect -228 942 -224 954
rect -210 946 -196 950
rect -172 948 -164 964
rect -159 957 -155 972
rect -144 954 -140 979
rect -113 973 -105 987
rect -100 965 -96 980
rect -105 961 -96 965
rect -124 954 -120 958
rect -100 955 -96 961
rect -144 950 -120 954
rect -54 954 -50 979
rect -23 973 -15 987
rect -10 965 -6 980
rect -15 961 -6 965
rect -34 954 -30 958
rect -10 955 -6 961
rect -54 950 -30 954
rect -144 948 -140 950
rect -172 944 -140 948
rect -172 942 -164 944
rect -188 938 -164 942
rect -203 905 -199 930
rect -172 924 -164 938
rect -54 941 -50 950
rect 18 941 22 1123
rect -54 937 22 941
rect 30 985 34 1123
rect 93 1136 97 1140
rect 93 1132 103 1136
rect 93 1120 97 1132
rect 111 1124 125 1128
rect 149 1126 157 1142
rect 162 1135 166 1150
rect 174 1126 178 1160
rect 205 1141 209 1160
rect 228 1157 232 1160
rect 252 1154 256 1160
rect 247 1150 256 1154
rect 149 1122 178 1126
rect 183 1136 187 1140
rect 183 1132 193 1136
rect 149 1120 157 1122
rect 183 1120 187 1132
rect 201 1124 215 1128
rect 239 1126 247 1142
rect 252 1135 256 1150
rect 239 1122 288 1126
rect 239 1120 247 1122
rect 133 1116 157 1120
rect 223 1116 247 1120
rect 118 1083 122 1108
rect 149 1102 157 1116
rect 162 1094 166 1109
rect 157 1090 166 1094
rect 138 1083 142 1087
rect 162 1084 166 1090
rect 118 1079 142 1083
rect 208 1083 212 1108
rect 239 1102 247 1116
rect 252 1094 256 1109
rect 247 1090 256 1094
rect 228 1083 232 1087
rect 252 1084 256 1090
rect 208 1079 232 1083
rect 118 1051 122 1079
rect 208 1070 212 1079
rect 208 1066 272 1070
rect 114 1047 123 1051
rect 119 1034 123 1047
rect 119 1030 146 1034
rect 178 1031 236 1034
rect 119 1011 123 1030
rect 142 1027 146 1030
rect 166 1024 170 1030
rect 161 1020 170 1024
rect 97 1006 101 1010
rect 97 1002 107 1006
rect 97 990 101 1002
rect 115 994 129 998
rect 153 996 161 1012
rect 166 1005 170 1020
rect 178 996 182 1031
rect 209 1030 236 1031
rect 209 1011 213 1030
rect 232 1027 236 1030
rect 256 1024 260 1030
rect 251 1020 260 1024
rect 153 992 182 996
rect 187 1006 191 1010
rect 187 1002 197 1006
rect 153 990 161 992
rect 187 990 191 1002
rect 205 994 219 998
rect 243 996 251 1012
rect 256 1005 260 1020
rect 268 996 272 1066
rect 243 992 272 996
rect 243 990 251 992
rect 137 986 161 990
rect 227 986 251 990
rect 30 981 87 985
rect -159 916 -155 931
rect -164 912 -155 916
rect -183 905 -179 909
rect -159 906 -155 912
rect -236 901 -179 905
rect 30 904 34 981
rect 60 962 64 981
rect 83 978 87 981
rect 107 975 111 981
rect 102 971 111 975
rect 38 957 42 961
rect 38 953 48 957
rect 38 941 42 953
rect 56 945 70 949
rect 94 947 102 963
rect 107 956 111 971
rect 122 953 126 978
rect 153 972 161 986
rect 166 964 170 979
rect 161 960 170 964
rect 142 953 146 957
rect 166 954 170 960
rect 122 949 146 953
rect 212 953 216 978
rect 243 972 251 986
rect 256 964 260 979
rect 251 960 260 964
rect 232 953 236 957
rect 256 954 260 960
rect 212 949 236 953
rect 122 947 126 949
rect 94 943 126 947
rect 94 941 102 943
rect 78 937 102 941
rect 63 904 67 929
rect 94 923 102 937
rect 212 940 216 949
rect 284 940 288 1122
rect 304 1000 308 1172
rect 328 1171 332 1172
rect 320 1158 324 1163
rect 316 1154 336 1158
rect 371 1153 375 1172
rect 394 1169 398 1172
rect 418 1166 422 1172
rect 413 1162 422 1166
rect 349 1148 353 1152
rect 349 1144 359 1148
rect 349 1132 353 1144
rect 367 1136 381 1140
rect 405 1138 413 1154
rect 418 1147 422 1162
rect 774 1156 798 1160
rect 987 1158 991 1333
rect 1072 1314 1076 1333
rect 1095 1330 1099 1333
rect 1119 1327 1123 1333
rect 1114 1323 1123 1327
rect 1050 1309 1054 1313
rect 1050 1305 1060 1309
rect 1050 1293 1054 1305
rect 1068 1297 1082 1301
rect 1106 1299 1114 1315
rect 1119 1308 1123 1323
rect 1131 1299 1135 1333
rect 1162 1314 1166 1333
rect 1185 1330 1189 1333
rect 1209 1327 1213 1333
rect 1204 1323 1213 1327
rect 1106 1295 1135 1299
rect 1140 1309 1144 1313
rect 1140 1305 1150 1309
rect 1106 1293 1114 1295
rect 1140 1293 1144 1305
rect 1158 1297 1172 1301
rect 1196 1299 1204 1315
rect 1209 1308 1213 1323
rect 1253 1332 1365 1336
rect 1397 1332 1455 1336
rect 1253 1299 1257 1332
rect 1338 1313 1342 1332
rect 1361 1329 1365 1332
rect 1385 1326 1389 1332
rect 1380 1322 1389 1326
rect 1196 1295 1257 1299
rect 1196 1293 1204 1295
rect 1090 1289 1114 1293
rect 1180 1289 1204 1293
rect 1075 1256 1079 1281
rect 1106 1275 1114 1289
rect 1119 1267 1123 1282
rect 1114 1263 1123 1267
rect 1095 1256 1099 1260
rect 1119 1257 1123 1263
rect 1075 1252 1099 1256
rect 1165 1256 1169 1281
rect 1196 1275 1204 1289
rect 1209 1267 1213 1282
rect 1204 1263 1213 1267
rect 1185 1256 1189 1260
rect 1209 1257 1213 1263
rect 1165 1252 1189 1256
rect 1035 1244 1059 1248
rect 1041 1239 1045 1244
rect 1049 1224 1053 1231
rect 1075 1224 1079 1252
rect 1165 1243 1169 1252
rect 1165 1239 1229 1243
rect 1030 1220 1034 1224
rect 1049 1220 1080 1224
rect 1049 1219 1053 1220
rect 1041 1206 1045 1211
rect 1076 1207 1080 1220
rect 1037 1202 1057 1206
rect 1076 1203 1103 1207
rect 1135 1204 1193 1207
rect 1076 1184 1080 1203
rect 1099 1200 1103 1203
rect 1123 1197 1127 1203
rect 1118 1193 1127 1197
rect 1054 1179 1058 1183
rect 1054 1175 1064 1179
rect 1054 1163 1058 1175
rect 1072 1167 1086 1171
rect 1110 1169 1118 1185
rect 1123 1178 1127 1193
rect 1135 1169 1139 1204
rect 1166 1203 1193 1204
rect 1166 1184 1170 1203
rect 1189 1200 1193 1203
rect 1213 1197 1217 1203
rect 1208 1193 1217 1197
rect 1110 1165 1139 1169
rect 1144 1179 1148 1183
rect 1144 1175 1154 1179
rect 1110 1163 1118 1165
rect 1144 1163 1148 1175
rect 1162 1167 1176 1171
rect 1200 1169 1208 1185
rect 1213 1178 1217 1193
rect 1225 1169 1229 1239
rect 1200 1165 1229 1169
rect 1200 1163 1208 1165
rect 1094 1159 1118 1163
rect 1184 1159 1208 1163
rect 780 1151 784 1156
rect 987 1154 1044 1158
rect 405 1134 461 1138
rect 788 1136 792 1143
rect 405 1132 413 1134
rect 389 1128 413 1132
rect 374 1109 378 1120
rect 405 1114 413 1128
rect 457 1131 461 1134
rect 764 1132 773 1136
rect 788 1132 858 1136
rect 457 1127 484 1131
rect 334 1105 378 1109
rect 418 1106 422 1121
rect 457 1108 461 1127
rect 480 1124 484 1127
rect 504 1121 508 1127
rect 499 1117 508 1121
rect 334 1101 338 1105
rect 316 1094 320 1098
rect 358 1094 362 1100
rect 316 1090 325 1094
rect 353 1090 362 1094
rect 374 1095 378 1105
rect 413 1102 422 1106
rect 394 1095 398 1099
rect 418 1096 422 1102
rect 435 1103 439 1107
rect 435 1099 445 1103
rect 374 1091 398 1095
rect 316 1078 320 1090
rect 333 1082 345 1086
rect 334 1071 338 1082
rect 358 1076 362 1090
rect 435 1087 439 1099
rect 453 1091 467 1095
rect 491 1093 499 1109
rect 504 1102 508 1117
rect 491 1089 514 1093
rect 491 1087 499 1089
rect 475 1083 499 1087
rect 371 1077 398 1081
rect 371 1071 375 1077
rect 334 1067 375 1071
rect 394 1074 398 1077
rect 418 1071 422 1077
rect 413 1067 422 1071
rect 371 1058 375 1067
rect 349 1053 353 1057
rect 349 1049 359 1053
rect 349 1037 353 1049
rect 367 1041 381 1045
rect 405 1043 413 1059
rect 418 1052 422 1067
rect 460 1050 464 1075
rect 491 1069 499 1083
rect 504 1061 508 1076
rect 499 1057 508 1061
rect 480 1050 484 1054
rect 504 1051 508 1057
rect 460 1046 484 1050
rect 527 1047 645 1051
rect 460 1043 464 1046
rect 405 1039 464 1043
rect 405 1037 413 1039
rect 389 1033 413 1037
rect 374 1000 378 1025
rect 405 1019 413 1033
rect 418 1011 422 1026
rect 527 1016 531 1047
rect 536 1036 560 1040
rect 542 1031 546 1036
rect 413 1007 422 1011
rect 394 1000 398 1004
rect 418 1001 422 1007
rect 513 1012 539 1016
rect 304 996 398 1000
rect 326 964 353 968
rect 326 945 330 964
rect 349 961 353 964
rect 373 958 377 964
rect 368 954 377 958
rect 212 936 288 940
rect 304 940 308 944
rect 304 936 314 940
rect 107 915 111 930
rect 304 924 308 936
rect 322 928 336 932
rect 360 930 368 946
rect 373 939 377 954
rect 391 950 415 954
rect 397 945 401 950
rect 405 930 409 937
rect 360 926 390 930
rect 405 926 426 930
rect 360 924 368 926
rect 405 925 409 926
rect 344 920 368 924
rect 102 911 111 915
rect 83 904 87 908
rect 107 905 111 911
rect 30 900 87 904
rect -236 889 -124 893
rect -92 889 -34 893
rect -236 714 -232 889
rect -151 870 -147 889
rect -128 886 -124 889
rect -104 883 -100 889
rect -109 879 -100 883
rect -173 865 -169 869
rect -173 861 -163 865
rect -173 849 -169 861
rect -155 853 -141 857
rect -117 855 -109 871
rect -104 864 -100 879
rect -92 855 -88 889
rect -61 870 -57 889
rect -38 886 -34 889
rect -14 883 -10 889
rect -19 879 -10 883
rect -117 851 -88 855
rect -83 865 -79 869
rect -83 861 -73 865
rect -117 849 -109 851
rect -83 849 -79 861
rect -65 853 -51 857
rect -27 855 -19 871
rect -14 864 -10 879
rect 30 888 142 892
rect 174 888 232 892
rect 30 855 34 888
rect 115 869 119 888
rect 138 885 142 888
rect 162 882 166 888
rect 157 878 166 882
rect -27 851 34 855
rect -27 849 -19 851
rect -133 845 -109 849
rect -43 845 -19 849
rect -148 812 -144 837
rect -117 831 -109 845
rect -104 823 -100 838
rect -109 819 -100 823
rect -128 812 -124 816
rect -104 813 -100 819
rect -148 808 -124 812
rect -58 812 -54 837
rect -27 831 -19 845
rect -14 823 -10 838
rect -19 819 -10 823
rect -38 812 -34 816
rect -14 813 -10 819
rect -58 808 -34 812
rect -188 800 -164 804
rect -182 795 -178 800
rect -174 780 -170 787
rect -148 780 -144 808
rect -58 799 -54 808
rect -58 795 6 799
rect -193 776 -189 780
rect -174 776 -143 780
rect -174 775 -170 776
rect -182 762 -178 767
rect -147 763 -143 776
rect -186 758 -166 762
rect -147 759 -120 763
rect -88 760 -30 763
rect -147 740 -143 759
rect -124 756 -120 759
rect -100 753 -96 759
rect -105 749 -96 753
rect -169 735 -165 739
rect -169 731 -159 735
rect -169 719 -165 731
rect -151 723 -137 727
rect -113 725 -105 741
rect -100 734 -96 749
rect -88 725 -84 760
rect -57 759 -30 760
rect -57 740 -53 759
rect -34 756 -30 759
rect -10 753 -6 759
rect -15 749 -6 753
rect -113 721 -84 725
rect -79 735 -75 739
rect -79 731 -69 735
rect -113 719 -105 721
rect -79 719 -75 731
rect -61 723 -47 727
rect -23 725 -15 741
rect -10 734 -6 749
rect 2 725 6 795
rect -23 721 6 725
rect -23 719 -15 721
rect -129 715 -105 719
rect -39 715 -15 719
rect -236 710 -179 714
rect -236 633 -232 710
rect -206 691 -202 710
rect -183 707 -179 710
rect -159 704 -155 710
rect -164 700 -155 704
rect -228 686 -224 690
rect -228 682 -218 686
rect -228 670 -224 682
rect -210 674 -196 678
rect -172 676 -164 692
rect -159 685 -155 700
rect -144 682 -140 707
rect -113 701 -105 715
rect -100 693 -96 708
rect -105 689 -96 693
rect -124 682 -120 686
rect -100 683 -96 689
rect -144 678 -120 682
rect -54 682 -50 707
rect -23 701 -15 715
rect -10 693 -6 708
rect -15 689 -6 693
rect -34 682 -30 686
rect -10 683 -6 689
rect -54 678 -30 682
rect -144 676 -140 678
rect -172 672 -140 676
rect -172 670 -164 672
rect -188 666 -164 670
rect -203 633 -199 658
rect -172 652 -164 666
rect -54 669 -50 678
rect 18 669 22 851
rect -54 665 22 669
rect 30 713 34 851
rect 93 864 97 868
rect 93 860 103 864
rect 93 848 97 860
rect 111 852 125 856
rect 149 854 157 870
rect 162 863 166 878
rect 174 854 178 888
rect 205 869 209 888
rect 228 885 232 888
rect 252 882 256 888
rect 329 887 333 912
rect 360 906 368 920
rect 373 898 377 913
rect 397 912 401 917
rect 393 908 413 912
rect 368 894 377 898
rect 349 887 353 891
rect 373 888 377 894
rect 329 883 353 887
rect 247 878 256 882
rect 149 850 178 854
rect 183 864 187 868
rect 183 860 193 864
rect 149 848 157 850
rect 183 848 187 860
rect 201 852 215 856
rect 239 854 247 870
rect 252 863 256 878
rect 314 861 338 865
rect 320 856 324 861
rect 239 850 288 854
rect 239 848 247 850
rect 133 844 157 848
rect 223 844 247 848
rect 118 811 122 836
rect 149 830 157 844
rect 162 822 166 837
rect 157 818 166 822
rect 138 811 142 815
rect 162 812 166 818
rect 118 807 142 811
rect 208 811 212 836
rect 239 830 247 844
rect 252 822 256 837
rect 247 818 256 822
rect 228 811 232 815
rect 252 812 256 818
rect 208 807 232 811
rect 118 779 122 807
rect 208 798 212 807
rect 208 794 272 798
rect 114 775 123 779
rect 119 762 123 775
rect 119 758 146 762
rect 178 759 236 762
rect 119 739 123 758
rect 142 755 146 758
rect 166 752 170 758
rect 161 748 170 752
rect 97 734 101 738
rect 97 730 107 734
rect 97 718 101 730
rect 115 722 129 726
rect 153 724 161 740
rect 166 733 170 748
rect 178 724 182 759
rect 209 758 236 759
rect 209 739 213 758
rect 232 755 236 758
rect 256 752 260 758
rect 251 748 260 752
rect 153 720 182 724
rect 187 734 191 738
rect 187 730 197 734
rect 153 718 161 720
rect 187 718 191 730
rect 205 722 219 726
rect 243 724 251 740
rect 256 733 260 748
rect 268 724 272 794
rect 243 720 272 724
rect 243 718 251 720
rect 137 714 161 718
rect 227 714 251 718
rect 30 709 87 713
rect -159 644 -155 659
rect -164 640 -155 644
rect -183 633 -179 637
rect -159 634 -155 640
rect -236 629 -179 633
rect 30 632 34 709
rect 60 690 64 709
rect 83 706 87 709
rect 107 703 111 709
rect 102 699 111 703
rect 38 685 42 689
rect 38 681 48 685
rect 38 669 42 681
rect 56 673 70 677
rect 94 675 102 691
rect 107 684 111 699
rect 122 681 126 706
rect 153 700 161 714
rect 166 692 170 707
rect 161 688 170 692
rect 142 681 146 685
rect 166 682 170 688
rect 122 677 146 681
rect 212 681 216 706
rect 243 700 251 714
rect 256 692 260 707
rect 251 688 260 692
rect 232 681 236 685
rect 256 682 260 688
rect 212 677 236 681
rect 122 675 126 677
rect 94 671 126 675
rect 94 669 102 671
rect 78 665 102 669
rect 63 632 67 657
rect 94 651 102 665
rect 212 668 216 677
rect 284 668 288 850
rect 328 841 332 848
rect 212 664 288 668
rect 304 837 313 841
rect 328 837 398 841
rect 304 665 308 837
rect 328 836 332 837
rect 320 823 324 828
rect 316 819 336 823
rect 371 818 375 837
rect 394 834 398 837
rect 418 831 422 837
rect 413 827 422 831
rect 349 813 353 817
rect 349 809 359 813
rect 349 797 353 809
rect 367 801 381 805
rect 405 803 413 819
rect 418 812 422 827
rect 513 818 517 1012
rect 550 897 554 1023
rect 565 1016 569 1047
rect 574 1036 598 1040
rect 580 1031 584 1036
rect 565 1012 577 1016
rect 588 938 592 1023
rect 603 1016 607 1047
rect 612 1036 636 1040
rect 618 1031 622 1036
rect 603 1012 615 1016
rect 626 979 630 1023
rect 641 1016 645 1047
rect 650 1036 674 1040
rect 719 1037 743 1041
rect 656 1031 660 1036
rect 725 1032 729 1037
rect 641 1012 653 1016
rect 664 1004 668 1023
rect 733 1017 737 1024
rect 712 1013 718 1017
rect 733 1013 748 1017
rect 733 1012 737 1013
rect 664 1000 698 1004
rect 664 991 668 1000
rect 694 992 698 1000
rect 725 999 729 1004
rect 721 995 741 999
rect 656 979 660 983
rect 626 975 660 979
rect 676 976 680 980
rect 626 950 630 975
rect 639 965 643 969
rect 656 961 660 975
rect 618 938 622 942
rect 588 934 622 938
rect 638 935 642 939
rect 588 909 592 934
rect 601 924 605 928
rect 618 920 622 934
rect 580 897 584 901
rect 550 893 584 897
rect 600 894 604 898
rect 533 872 537 876
rect 550 868 554 893
rect 563 883 567 887
rect 580 879 584 893
rect 525 843 529 847
rect 542 839 546 860
rect 534 821 538 831
rect 572 821 576 871
rect 610 821 614 912
rect 648 821 652 953
rect 686 821 690 984
rect 706 977 710 981
rect 719 980 743 984
rect 725 975 729 980
rect 733 960 737 967
rect 764 960 768 1132
rect 788 1131 792 1132
rect 780 1118 784 1123
rect 776 1114 796 1118
rect 831 1113 835 1132
rect 854 1129 858 1132
rect 878 1126 882 1132
rect 873 1122 882 1126
rect 809 1108 813 1112
rect 809 1104 819 1108
rect 809 1092 813 1104
rect 827 1096 841 1100
rect 865 1098 873 1114
rect 878 1107 882 1122
rect 865 1094 921 1098
rect 865 1092 873 1094
rect 849 1088 873 1092
rect 834 1069 838 1080
rect 865 1074 873 1088
rect 917 1091 921 1094
rect 917 1087 944 1091
rect 794 1065 838 1069
rect 878 1066 882 1081
rect 917 1068 921 1087
rect 940 1084 944 1087
rect 964 1081 968 1087
rect 959 1077 968 1081
rect 794 1061 798 1065
rect 776 1054 780 1058
rect 818 1054 822 1060
rect 776 1050 785 1054
rect 813 1050 822 1054
rect 834 1055 838 1065
rect 873 1062 882 1066
rect 854 1055 858 1059
rect 878 1056 882 1062
rect 895 1063 899 1067
rect 895 1059 905 1063
rect 834 1051 858 1055
rect 776 1038 780 1050
rect 793 1042 805 1046
rect 794 1031 798 1042
rect 818 1036 822 1050
rect 895 1047 899 1059
rect 913 1051 927 1055
rect 951 1053 959 1069
rect 964 1062 968 1077
rect 987 1077 991 1154
rect 1017 1135 1021 1154
rect 1040 1151 1044 1154
rect 1064 1148 1068 1154
rect 1059 1144 1068 1148
rect 995 1130 999 1134
rect 995 1126 1005 1130
rect 995 1114 999 1126
rect 1013 1118 1027 1122
rect 1051 1120 1059 1136
rect 1064 1129 1068 1144
rect 1079 1126 1083 1151
rect 1110 1145 1118 1159
rect 1123 1137 1127 1152
rect 1118 1133 1127 1137
rect 1099 1126 1103 1130
rect 1123 1127 1127 1133
rect 1079 1122 1103 1126
rect 1169 1126 1173 1151
rect 1200 1145 1208 1159
rect 1213 1137 1217 1152
rect 1208 1133 1217 1137
rect 1189 1126 1193 1130
rect 1213 1127 1217 1133
rect 1169 1122 1193 1126
rect 1079 1120 1083 1122
rect 1051 1116 1083 1120
rect 1051 1114 1059 1116
rect 1035 1110 1059 1114
rect 1020 1077 1024 1102
rect 1051 1096 1059 1110
rect 1169 1113 1173 1122
rect 1241 1113 1245 1295
rect 1169 1109 1245 1113
rect 1253 1157 1257 1295
rect 1316 1308 1320 1312
rect 1316 1304 1326 1308
rect 1316 1292 1320 1304
rect 1334 1296 1348 1300
rect 1372 1298 1380 1314
rect 1385 1307 1389 1322
rect 1397 1298 1401 1332
rect 1428 1313 1432 1332
rect 1451 1329 1455 1332
rect 1475 1326 1479 1332
rect 1470 1322 1479 1326
rect 1372 1294 1401 1298
rect 1406 1308 1410 1312
rect 1406 1304 1416 1308
rect 1372 1292 1380 1294
rect 1406 1292 1410 1304
rect 1424 1296 1438 1300
rect 1462 1298 1470 1314
rect 1475 1307 1479 1322
rect 1462 1294 1511 1298
rect 1462 1292 1470 1294
rect 1356 1288 1380 1292
rect 1446 1288 1470 1292
rect 1341 1255 1345 1280
rect 1372 1274 1380 1288
rect 1385 1266 1389 1281
rect 1380 1262 1389 1266
rect 1361 1255 1365 1259
rect 1385 1256 1389 1262
rect 1341 1251 1365 1255
rect 1431 1255 1435 1280
rect 1462 1274 1470 1288
rect 1475 1266 1479 1281
rect 1470 1262 1479 1266
rect 1451 1255 1455 1259
rect 1475 1256 1479 1262
rect 1431 1251 1455 1255
rect 1341 1223 1345 1251
rect 1431 1242 1435 1251
rect 1431 1238 1495 1242
rect 1337 1219 1346 1223
rect 1342 1206 1346 1219
rect 1342 1202 1369 1206
rect 1401 1203 1459 1206
rect 1342 1183 1346 1202
rect 1365 1199 1369 1202
rect 1389 1196 1393 1202
rect 1384 1192 1393 1196
rect 1320 1178 1324 1182
rect 1320 1174 1330 1178
rect 1320 1162 1324 1174
rect 1338 1166 1352 1170
rect 1376 1168 1384 1184
rect 1389 1177 1393 1192
rect 1401 1168 1405 1203
rect 1432 1202 1459 1203
rect 1432 1183 1436 1202
rect 1455 1199 1459 1202
rect 1479 1196 1483 1202
rect 1474 1192 1483 1196
rect 1376 1164 1405 1168
rect 1410 1178 1414 1182
rect 1410 1174 1420 1178
rect 1376 1162 1384 1164
rect 1410 1162 1414 1174
rect 1428 1166 1442 1170
rect 1466 1168 1474 1184
rect 1479 1177 1483 1192
rect 1491 1168 1495 1238
rect 1466 1164 1495 1168
rect 1466 1162 1474 1164
rect 1360 1158 1384 1162
rect 1450 1158 1474 1162
rect 1253 1153 1310 1157
rect 1064 1088 1068 1103
rect 1059 1084 1068 1088
rect 1040 1077 1044 1081
rect 1064 1078 1068 1084
rect 987 1073 1044 1077
rect 1253 1076 1257 1153
rect 1283 1134 1287 1153
rect 1306 1150 1310 1153
rect 1330 1147 1334 1153
rect 1325 1143 1334 1147
rect 1261 1129 1265 1133
rect 1261 1125 1271 1129
rect 1261 1113 1265 1125
rect 1279 1117 1293 1121
rect 1317 1119 1325 1135
rect 1330 1128 1334 1143
rect 1345 1125 1349 1150
rect 1376 1144 1384 1158
rect 1389 1136 1393 1151
rect 1384 1132 1393 1136
rect 1365 1125 1369 1129
rect 1389 1126 1393 1132
rect 1345 1121 1369 1125
rect 1435 1125 1439 1150
rect 1466 1144 1474 1158
rect 1479 1136 1483 1151
rect 1474 1132 1483 1136
rect 1455 1125 1459 1129
rect 1479 1126 1483 1132
rect 1435 1121 1459 1125
rect 1345 1119 1349 1121
rect 1317 1115 1349 1119
rect 1317 1113 1325 1115
rect 1301 1109 1325 1113
rect 1286 1076 1290 1101
rect 1317 1095 1325 1109
rect 1435 1112 1439 1121
rect 1507 1112 1511 1294
rect 1435 1108 1511 1112
rect 1330 1087 1334 1102
rect 1325 1083 1334 1087
rect 1306 1076 1310 1080
rect 1330 1077 1334 1083
rect 1253 1072 1310 1076
rect 987 1061 1099 1065
rect 1131 1061 1189 1065
rect 951 1049 971 1053
rect 951 1047 959 1049
rect 935 1043 959 1047
rect 831 1037 858 1041
rect 831 1031 835 1037
rect 794 1027 835 1031
rect 854 1034 858 1037
rect 878 1031 882 1037
rect 873 1027 882 1031
rect 831 1018 835 1027
rect 809 1013 813 1017
rect 809 1009 819 1013
rect 809 997 813 1009
rect 827 1001 841 1005
rect 865 1003 873 1019
rect 878 1012 882 1027
rect 920 1010 924 1035
rect 951 1029 959 1043
rect 964 1021 968 1036
rect 959 1017 968 1021
rect 940 1010 944 1014
rect 964 1011 968 1017
rect 920 1006 944 1010
rect 920 1003 924 1006
rect 865 999 924 1003
rect 865 997 873 999
rect 849 993 873 997
rect 834 960 838 985
rect 865 979 873 993
rect 878 971 882 986
rect 873 967 882 971
rect 854 960 858 964
rect 878 961 882 967
rect 712 956 718 960
rect 733 956 748 960
rect 764 956 858 960
rect 733 955 737 956
rect 725 942 729 947
rect 721 938 741 942
rect 719 923 743 927
rect 774 923 798 927
rect 725 918 729 923
rect 780 918 784 923
rect 733 903 737 910
rect 788 903 792 910
rect 712 899 718 903
rect 733 899 748 903
rect 764 899 773 903
rect 788 899 858 903
rect 733 898 737 899
rect 725 885 729 890
rect 721 881 741 885
rect 719 866 743 870
rect 725 861 729 866
rect 733 846 737 853
rect 712 842 718 846
rect 733 842 748 846
rect 733 841 737 842
rect 725 828 729 833
rect 721 824 741 828
rect 513 814 521 818
rect 534 817 690 821
rect 534 810 538 817
rect 405 799 461 803
rect 405 797 413 799
rect 389 793 413 797
rect 374 774 378 785
rect 405 779 413 793
rect 457 796 461 799
rect 526 796 530 802
rect 457 792 484 796
rect 522 792 542 796
rect 334 770 378 774
rect 418 771 422 786
rect 457 773 461 792
rect 480 789 484 792
rect 504 786 508 792
rect 499 782 508 786
rect 334 766 338 770
rect 316 759 320 763
rect 358 759 362 765
rect 316 755 325 759
rect 353 755 362 759
rect 374 760 378 770
rect 413 767 422 771
rect 394 760 398 764
rect 418 761 422 767
rect 435 768 439 772
rect 435 764 445 768
rect 374 756 398 760
rect 316 743 320 755
rect 333 747 345 751
rect 334 736 338 747
rect 358 741 362 755
rect 435 752 439 764
rect 453 756 467 760
rect 491 758 499 774
rect 504 767 508 782
rect 491 754 514 758
rect 491 752 499 754
rect 475 748 499 752
rect 371 742 398 746
rect 371 736 375 742
rect 334 732 375 736
rect 394 739 398 742
rect 418 736 422 742
rect 413 732 422 736
rect 371 723 375 732
rect 349 718 353 722
rect 349 714 359 718
rect 349 702 353 714
rect 367 706 381 710
rect 405 708 413 724
rect 418 717 422 732
rect 460 715 464 740
rect 491 734 499 748
rect 504 726 508 741
rect 499 722 508 726
rect 764 727 768 899
rect 788 898 792 899
rect 780 885 784 890
rect 776 881 796 885
rect 831 880 835 899
rect 854 896 858 899
rect 878 893 882 899
rect 873 889 882 893
rect 809 875 813 879
rect 809 871 819 875
rect 809 859 813 871
rect 827 863 841 867
rect 865 865 873 881
rect 878 874 882 889
rect 987 886 991 1061
rect 1072 1042 1076 1061
rect 1095 1058 1099 1061
rect 1119 1055 1123 1061
rect 1114 1051 1123 1055
rect 1050 1037 1054 1041
rect 1050 1033 1060 1037
rect 1050 1021 1054 1033
rect 1068 1025 1082 1029
rect 1106 1027 1114 1043
rect 1119 1036 1123 1051
rect 1131 1027 1135 1061
rect 1162 1042 1166 1061
rect 1185 1058 1189 1061
rect 1209 1055 1213 1061
rect 1204 1051 1213 1055
rect 1106 1023 1135 1027
rect 1140 1037 1144 1041
rect 1140 1033 1150 1037
rect 1106 1021 1114 1023
rect 1140 1021 1144 1033
rect 1158 1025 1172 1029
rect 1196 1027 1204 1043
rect 1209 1036 1213 1051
rect 1253 1060 1365 1064
rect 1397 1060 1455 1064
rect 1253 1027 1257 1060
rect 1338 1041 1342 1060
rect 1361 1057 1365 1060
rect 1385 1054 1389 1060
rect 1380 1050 1389 1054
rect 1196 1023 1257 1027
rect 1196 1021 1204 1023
rect 1090 1017 1114 1021
rect 1180 1017 1204 1021
rect 1075 984 1079 1009
rect 1106 1003 1114 1017
rect 1119 995 1123 1010
rect 1114 991 1123 995
rect 1095 984 1099 988
rect 1119 985 1123 991
rect 1075 980 1099 984
rect 1165 984 1169 1009
rect 1196 1003 1204 1017
rect 1209 995 1213 1010
rect 1204 991 1213 995
rect 1185 984 1189 988
rect 1209 985 1213 991
rect 1165 980 1189 984
rect 1035 972 1059 976
rect 1041 967 1045 972
rect 1049 952 1053 959
rect 1075 952 1079 980
rect 1165 971 1169 980
rect 1165 967 1229 971
rect 1030 948 1034 952
rect 1049 948 1080 952
rect 1049 947 1053 948
rect 1041 934 1045 939
rect 1076 935 1080 948
rect 1037 930 1057 934
rect 1076 931 1103 935
rect 1135 932 1193 935
rect 1076 912 1080 931
rect 1099 928 1103 931
rect 1123 925 1127 931
rect 1118 921 1127 925
rect 1054 907 1058 911
rect 1054 903 1064 907
rect 1054 891 1058 903
rect 1072 895 1086 899
rect 1110 897 1118 913
rect 1123 906 1127 921
rect 1135 897 1139 932
rect 1166 931 1193 932
rect 1166 912 1170 931
rect 1189 928 1193 931
rect 1213 925 1217 931
rect 1208 921 1217 925
rect 1110 893 1139 897
rect 1144 907 1148 911
rect 1144 903 1154 907
rect 1110 891 1118 893
rect 1144 891 1148 903
rect 1162 895 1176 899
rect 1200 897 1208 913
rect 1213 906 1217 921
rect 1225 897 1229 967
rect 1200 893 1229 897
rect 1200 891 1208 893
rect 1094 887 1118 891
rect 1184 887 1208 891
rect 987 882 1044 886
rect 865 861 921 865
rect 865 859 873 861
rect 849 855 873 859
rect 834 836 838 847
rect 865 841 873 855
rect 917 858 921 861
rect 917 854 944 858
rect 794 832 838 836
rect 878 833 882 848
rect 917 835 921 854
rect 940 851 944 854
rect 964 848 968 854
rect 959 844 968 848
rect 794 828 798 832
rect 776 821 780 825
rect 818 821 822 827
rect 776 817 785 821
rect 813 817 822 821
rect 834 822 838 832
rect 873 829 882 833
rect 854 822 858 826
rect 878 823 882 829
rect 895 830 899 834
rect 895 826 905 830
rect 834 818 858 822
rect 776 805 780 817
rect 793 809 805 813
rect 794 798 798 809
rect 818 803 822 817
rect 895 814 899 826
rect 913 818 927 822
rect 951 820 959 836
rect 964 829 968 844
rect 951 816 971 820
rect 951 814 959 816
rect 935 810 959 814
rect 831 804 858 808
rect 831 798 835 804
rect 794 794 835 798
rect 854 801 858 804
rect 878 798 882 804
rect 873 794 882 798
rect 831 785 835 794
rect 809 780 813 784
rect 809 776 819 780
rect 809 764 813 776
rect 827 768 841 772
rect 865 770 873 786
rect 878 779 882 794
rect 920 777 924 802
rect 951 796 959 810
rect 987 805 991 882
rect 1017 863 1021 882
rect 1040 879 1044 882
rect 1064 876 1068 882
rect 1059 872 1068 876
rect 995 858 999 862
rect 995 854 1005 858
rect 995 842 999 854
rect 1013 846 1027 850
rect 1051 848 1059 864
rect 1064 857 1068 872
rect 1079 854 1083 879
rect 1110 873 1118 887
rect 1123 865 1127 880
rect 1118 861 1127 865
rect 1099 854 1103 858
rect 1123 855 1127 861
rect 1079 850 1103 854
rect 1169 854 1173 879
rect 1200 873 1208 887
rect 1213 865 1217 880
rect 1208 861 1217 865
rect 1189 854 1193 858
rect 1213 855 1217 861
rect 1169 850 1193 854
rect 1079 848 1083 850
rect 1051 844 1083 848
rect 1051 842 1059 844
rect 1035 838 1059 842
rect 1020 805 1024 830
rect 1051 824 1059 838
rect 1169 841 1173 850
rect 1241 841 1245 1023
rect 1169 837 1245 841
rect 1253 885 1257 1023
rect 1316 1036 1320 1040
rect 1316 1032 1326 1036
rect 1316 1020 1320 1032
rect 1334 1024 1348 1028
rect 1372 1026 1380 1042
rect 1385 1035 1389 1050
rect 1397 1026 1401 1060
rect 1428 1041 1432 1060
rect 1451 1057 1455 1060
rect 1475 1054 1479 1060
rect 1470 1050 1479 1054
rect 1372 1022 1401 1026
rect 1406 1036 1410 1040
rect 1406 1032 1416 1036
rect 1372 1020 1380 1022
rect 1406 1020 1410 1032
rect 1424 1024 1438 1028
rect 1462 1026 1470 1042
rect 1475 1035 1479 1050
rect 1462 1022 1511 1026
rect 1462 1020 1470 1022
rect 1356 1016 1380 1020
rect 1446 1016 1470 1020
rect 1341 983 1345 1008
rect 1372 1002 1380 1016
rect 1385 994 1389 1009
rect 1380 990 1389 994
rect 1361 983 1365 987
rect 1385 984 1389 990
rect 1341 979 1365 983
rect 1431 983 1435 1008
rect 1462 1002 1470 1016
rect 1475 994 1479 1009
rect 1470 990 1479 994
rect 1451 983 1455 987
rect 1475 984 1479 990
rect 1431 979 1455 983
rect 1341 951 1345 979
rect 1431 970 1435 979
rect 1431 966 1495 970
rect 1337 947 1346 951
rect 1342 934 1346 947
rect 1342 930 1369 934
rect 1401 931 1459 934
rect 1342 911 1346 930
rect 1365 927 1369 930
rect 1389 924 1393 930
rect 1384 920 1393 924
rect 1320 906 1324 910
rect 1320 902 1330 906
rect 1320 890 1324 902
rect 1338 894 1352 898
rect 1376 896 1384 912
rect 1389 905 1393 920
rect 1401 896 1405 931
rect 1432 930 1459 931
rect 1432 911 1436 930
rect 1455 927 1459 930
rect 1479 924 1483 930
rect 1474 920 1483 924
rect 1376 892 1405 896
rect 1410 906 1414 910
rect 1410 902 1420 906
rect 1376 890 1384 892
rect 1410 890 1414 902
rect 1428 894 1442 898
rect 1466 896 1474 912
rect 1479 905 1483 920
rect 1491 896 1495 966
rect 1466 892 1495 896
rect 1466 890 1474 892
rect 1360 886 1384 890
rect 1450 886 1474 890
rect 1253 881 1310 885
rect 1064 816 1068 831
rect 1059 812 1068 816
rect 1040 805 1044 809
rect 1064 806 1068 812
rect 964 788 968 803
rect 987 801 1044 805
rect 1253 804 1257 881
rect 1283 862 1287 881
rect 1306 878 1310 881
rect 1330 875 1334 881
rect 1325 871 1334 875
rect 1261 857 1265 861
rect 1261 853 1271 857
rect 1261 841 1265 853
rect 1279 845 1293 849
rect 1317 847 1325 863
rect 1330 856 1334 871
rect 1345 853 1349 878
rect 1376 872 1384 886
rect 1389 864 1393 879
rect 1384 860 1393 864
rect 1365 853 1369 857
rect 1389 854 1393 860
rect 1345 849 1369 853
rect 1435 853 1439 878
rect 1466 872 1474 886
rect 1479 864 1483 879
rect 1474 860 1483 864
rect 1455 853 1459 857
rect 1479 854 1483 860
rect 1435 849 1459 853
rect 1345 847 1349 849
rect 1317 843 1349 847
rect 1317 841 1325 843
rect 1301 837 1325 841
rect 1286 804 1290 829
rect 1317 823 1325 837
rect 1435 840 1439 849
rect 1507 840 1511 1022
rect 1435 836 1511 840
rect 1330 815 1334 830
rect 1325 811 1334 815
rect 1306 804 1310 808
rect 1330 805 1334 811
rect 1253 800 1310 804
rect 959 784 968 788
rect 940 777 944 781
rect 964 778 968 784
rect 987 789 1099 793
rect 1131 789 1189 793
rect 920 773 944 777
rect 920 770 924 773
rect 865 766 924 770
rect 865 764 873 766
rect 849 760 873 764
rect 834 727 838 752
rect 865 746 873 760
rect 878 738 882 753
rect 873 734 882 738
rect 854 727 858 731
rect 878 728 882 734
rect 764 723 858 727
rect 480 715 484 719
rect 504 716 508 722
rect 460 711 484 715
rect 460 708 464 711
rect 405 704 464 708
rect 405 702 413 704
rect 389 698 413 702
rect 374 665 378 690
rect 405 684 413 698
rect 418 676 422 691
rect 774 690 798 694
rect 780 685 784 690
rect 413 672 422 676
rect 394 665 398 669
rect 418 666 422 672
rect 788 670 792 677
rect 764 666 773 670
rect 788 666 858 670
rect 304 661 398 665
rect 107 643 111 658
rect 102 639 111 643
rect 83 632 87 636
rect 107 633 111 639
rect 30 628 87 632
rect 326 629 353 633
rect -236 617 -124 621
rect -92 617 -34 621
rect -236 442 -232 617
rect -151 598 -147 617
rect -128 614 -124 617
rect -104 611 -100 617
rect -109 607 -100 611
rect -173 593 -169 597
rect -173 589 -163 593
rect -173 577 -169 589
rect -155 581 -141 585
rect -117 583 -109 599
rect -104 592 -100 607
rect -92 583 -88 617
rect -61 598 -57 617
rect -38 614 -34 617
rect -14 611 -10 617
rect -19 607 -10 611
rect -117 579 -88 583
rect -83 593 -79 597
rect -83 589 -73 593
rect -117 577 -109 579
rect -83 577 -79 589
rect -65 581 -51 585
rect -27 583 -19 599
rect -14 592 -10 607
rect 30 616 142 620
rect 174 616 232 620
rect 30 583 34 616
rect 115 597 119 616
rect 138 613 142 616
rect 162 610 166 616
rect 157 606 166 610
rect -27 579 34 583
rect -27 577 -19 579
rect -133 573 -109 577
rect -43 573 -19 577
rect -148 540 -144 565
rect -117 559 -109 573
rect -104 551 -100 566
rect -109 547 -100 551
rect -128 540 -124 544
rect -104 541 -100 547
rect -148 536 -124 540
rect -58 540 -54 565
rect -27 559 -19 573
rect -14 551 -10 566
rect -19 547 -10 551
rect -38 540 -34 544
rect -14 541 -10 547
rect -58 536 -34 540
rect -188 528 -164 532
rect -182 523 -178 528
rect -174 508 -170 515
rect -148 508 -144 536
rect -58 527 -54 536
rect -58 523 6 527
rect -193 504 -189 508
rect -174 504 -143 508
rect -174 503 -170 504
rect -182 490 -178 495
rect -147 491 -143 504
rect -186 486 -166 490
rect -147 487 -120 491
rect -88 488 -30 491
rect -147 468 -143 487
rect -124 484 -120 487
rect -100 481 -96 487
rect -105 477 -96 481
rect -169 463 -165 467
rect -169 459 -159 463
rect -169 447 -165 459
rect -151 451 -137 455
rect -113 453 -105 469
rect -100 462 -96 477
rect -88 453 -84 488
rect -57 487 -30 488
rect -57 468 -53 487
rect -34 484 -30 487
rect -10 481 -6 487
rect -15 477 -6 481
rect -113 449 -84 453
rect -79 463 -75 467
rect -79 459 -69 463
rect -113 447 -105 449
rect -79 447 -75 459
rect -61 451 -47 455
rect -23 453 -15 469
rect -10 462 -6 477
rect 2 453 6 523
rect -23 449 6 453
rect -23 447 -15 449
rect -129 443 -105 447
rect -39 443 -15 447
rect -236 438 -179 442
rect -236 361 -232 438
rect -206 419 -202 438
rect -183 435 -179 438
rect -159 432 -155 438
rect -164 428 -155 432
rect -228 414 -224 418
rect -228 410 -218 414
rect -228 398 -224 410
rect -210 402 -196 406
rect -172 404 -164 420
rect -159 413 -155 428
rect -144 410 -140 435
rect -113 429 -105 443
rect -100 421 -96 436
rect -105 417 -96 421
rect -124 410 -120 414
rect -100 411 -96 417
rect -144 406 -120 410
rect -54 410 -50 435
rect -23 429 -15 443
rect -10 421 -6 436
rect -15 417 -6 421
rect -34 410 -30 414
rect -10 411 -6 417
rect -54 406 -30 410
rect -144 404 -140 406
rect -172 400 -140 404
rect -172 398 -164 400
rect -188 394 -164 398
rect -203 361 -199 386
rect -172 380 -164 394
rect -54 397 -50 406
rect 18 397 22 579
rect -54 393 22 397
rect 30 441 34 579
rect 93 592 97 596
rect 93 588 103 592
rect 93 576 97 588
rect 111 580 125 584
rect 149 582 157 598
rect 162 591 166 606
rect 174 582 178 616
rect 205 597 209 616
rect 228 613 232 616
rect 252 610 256 616
rect 247 606 256 610
rect 326 610 330 629
rect 349 626 353 629
rect 373 623 377 629
rect 368 619 377 623
rect 149 578 178 582
rect 183 592 187 596
rect 183 588 193 592
rect 149 576 157 578
rect 183 576 187 588
rect 201 580 215 584
rect 239 582 247 598
rect 252 591 256 606
rect 304 605 308 609
rect 304 601 314 605
rect 304 589 308 601
rect 322 593 336 597
rect 360 595 368 611
rect 373 604 377 619
rect 391 615 415 619
rect 397 610 401 615
rect 405 595 409 602
rect 360 591 390 595
rect 405 591 426 595
rect 360 589 368 591
rect 405 590 409 591
rect 344 585 368 589
rect 239 578 288 582
rect 239 576 247 578
rect 133 572 157 576
rect 223 572 247 576
rect 118 539 122 564
rect 149 558 157 572
rect 162 550 166 565
rect 157 546 166 550
rect 138 539 142 543
rect 162 540 166 546
rect 118 535 142 539
rect 208 539 212 564
rect 239 558 247 572
rect 252 550 256 565
rect 247 546 256 550
rect 228 539 232 543
rect 252 540 256 546
rect 208 535 232 539
rect 118 507 122 535
rect 208 526 212 535
rect 208 522 272 526
rect 114 503 123 507
rect 119 490 123 503
rect 119 486 146 490
rect 178 487 236 490
rect 119 467 123 486
rect 142 483 146 486
rect 166 480 170 486
rect 161 476 170 480
rect 97 462 101 466
rect 97 458 107 462
rect 97 446 101 458
rect 115 450 129 454
rect 153 452 161 468
rect 166 461 170 476
rect 178 452 182 487
rect 209 486 236 487
rect 209 467 213 486
rect 232 483 236 486
rect 256 480 260 486
rect 251 476 260 480
rect 153 448 182 452
rect 187 462 191 466
rect 187 458 197 462
rect 153 446 161 448
rect 187 446 191 458
rect 205 450 219 454
rect 243 452 251 468
rect 256 461 260 476
rect 268 452 272 522
rect 243 448 272 452
rect 243 446 251 448
rect 137 442 161 446
rect 227 442 251 446
rect 30 437 87 441
rect -159 372 -155 387
rect -164 368 -155 372
rect -183 361 -179 365
rect -159 362 -155 368
rect -236 357 -179 361
rect 30 360 34 437
rect 60 418 64 437
rect 83 434 87 437
rect 107 431 111 437
rect 102 427 111 431
rect 38 413 42 417
rect 38 409 48 413
rect 38 397 42 409
rect 56 401 70 405
rect 94 403 102 419
rect 107 412 111 427
rect 122 409 126 434
rect 153 428 161 442
rect 166 420 170 435
rect 161 416 170 420
rect 142 409 146 413
rect 166 410 170 416
rect 122 405 146 409
rect 212 409 216 434
rect 243 428 251 442
rect 256 420 260 435
rect 251 416 260 420
rect 232 409 236 413
rect 256 410 260 416
rect 212 405 236 409
rect 122 403 126 405
rect 94 399 126 403
rect 94 397 102 399
rect 78 393 102 397
rect 63 360 67 385
rect 94 379 102 393
rect 212 396 216 405
rect 284 396 288 578
rect 329 552 333 577
rect 360 571 368 585
rect 373 563 377 578
rect 397 577 401 582
rect 393 573 413 577
rect 368 559 377 563
rect 349 552 353 556
rect 373 553 377 559
rect 329 548 353 552
rect 314 526 338 530
rect 320 521 324 526
rect 328 506 332 513
rect 212 392 288 396
rect 304 502 313 506
rect 328 502 398 506
rect 107 371 111 386
rect 102 367 111 371
rect 83 360 87 364
rect 107 361 111 367
rect 30 356 87 360
rect -236 345 -124 349
rect -92 345 -34 349
rect -236 170 -232 345
rect -151 326 -147 345
rect -128 342 -124 345
rect -104 339 -100 345
rect -109 335 -100 339
rect -173 321 -169 325
rect -173 317 -163 321
rect -173 305 -169 317
rect -155 309 -141 313
rect -117 311 -109 327
rect -104 320 -100 335
rect -92 311 -88 345
rect -61 326 -57 345
rect -38 342 -34 345
rect -14 339 -10 345
rect -19 335 -10 339
rect -117 307 -88 311
rect -83 321 -79 325
rect -83 317 -73 321
rect -117 305 -109 307
rect -83 305 -79 317
rect -65 309 -51 313
rect -27 311 -19 327
rect -14 320 -10 335
rect 30 344 142 348
rect 174 344 232 348
rect 30 311 34 344
rect 115 325 119 344
rect 138 341 142 344
rect 162 338 166 344
rect 157 334 166 338
rect -27 307 34 311
rect -27 305 -19 307
rect -133 301 -109 305
rect -43 301 -19 305
rect -148 268 -144 293
rect -117 287 -109 301
rect -104 279 -100 294
rect -109 275 -100 279
rect -128 268 -124 272
rect -104 269 -100 275
rect -148 264 -124 268
rect -58 268 -54 293
rect -27 287 -19 301
rect -14 279 -10 294
rect -19 275 -10 279
rect -38 268 -34 272
rect -14 269 -10 275
rect -58 264 -34 268
rect -188 256 -164 260
rect -182 251 -178 256
rect -174 236 -170 243
rect -148 236 -144 264
rect -58 255 -54 264
rect -58 251 6 255
rect -193 232 -189 236
rect -174 232 -143 236
rect -174 231 -170 232
rect -182 218 -178 223
rect -147 219 -143 232
rect -186 214 -166 218
rect -147 215 -120 219
rect -88 216 -30 219
rect -147 196 -143 215
rect -124 212 -120 215
rect -100 209 -96 215
rect -105 205 -96 209
rect -169 191 -165 195
rect -169 187 -159 191
rect -169 175 -165 187
rect -151 179 -137 183
rect -113 181 -105 197
rect -100 190 -96 205
rect -88 181 -84 216
rect -57 215 -30 216
rect -57 196 -53 215
rect -34 212 -30 215
rect -10 209 -6 215
rect -15 205 -6 209
rect -113 177 -84 181
rect -79 191 -75 195
rect -79 187 -69 191
rect -113 175 -105 177
rect -79 175 -75 187
rect -61 179 -47 183
rect -23 181 -15 197
rect -10 190 -6 205
rect 2 181 6 251
rect -23 177 6 181
rect -23 175 -15 177
rect -129 171 -105 175
rect -39 171 -15 175
rect -236 166 -179 170
rect -236 89 -232 166
rect -206 147 -202 166
rect -183 163 -179 166
rect -159 160 -155 166
rect -164 156 -155 160
rect -228 142 -224 146
rect -228 138 -218 142
rect -228 126 -224 138
rect -210 130 -196 134
rect -172 132 -164 148
rect -159 141 -155 156
rect -144 138 -140 163
rect -113 157 -105 171
rect -100 149 -96 164
rect -105 145 -96 149
rect -124 138 -120 142
rect -100 139 -96 145
rect -144 134 -120 138
rect -54 138 -50 163
rect -23 157 -15 171
rect -10 149 -6 164
rect -15 145 -6 149
rect -34 138 -30 142
rect -10 139 -6 145
rect -54 134 -30 138
rect -144 132 -140 134
rect -172 128 -140 132
rect -172 126 -164 128
rect -188 122 -164 126
rect -203 89 -199 114
rect -172 108 -164 122
rect -54 125 -50 134
rect 18 125 22 307
rect -54 121 22 125
rect 30 169 34 307
rect 93 320 97 324
rect 93 316 103 320
rect 93 304 97 316
rect 111 308 125 312
rect 149 310 157 326
rect 162 319 166 334
rect 174 310 178 344
rect 205 325 209 344
rect 228 341 232 344
rect 252 338 256 344
rect 247 334 256 338
rect 149 306 178 310
rect 183 320 187 324
rect 183 316 193 320
rect 149 304 157 306
rect 183 304 187 316
rect 201 308 215 312
rect 239 310 247 326
rect 252 319 256 334
rect 304 330 308 502
rect 328 501 332 502
rect 320 488 324 493
rect 316 484 336 488
rect 371 483 375 502
rect 394 499 398 502
rect 418 496 422 502
rect 413 492 422 496
rect 349 478 353 482
rect 349 474 359 478
rect 349 462 353 474
rect 367 466 381 470
rect 405 468 413 484
rect 418 477 422 492
rect 764 494 768 666
rect 788 665 792 666
rect 780 652 784 657
rect 776 648 796 652
rect 831 647 835 666
rect 854 663 858 666
rect 878 660 882 666
rect 873 656 882 660
rect 809 642 813 646
rect 809 638 819 642
rect 809 626 813 638
rect 827 630 841 634
rect 865 632 873 648
rect 878 641 882 656
rect 865 628 921 632
rect 865 626 873 628
rect 849 622 873 626
rect 834 603 838 614
rect 865 608 873 622
rect 917 625 921 628
rect 917 621 944 625
rect 794 599 838 603
rect 878 600 882 615
rect 917 602 921 621
rect 940 618 944 621
rect 964 615 968 621
rect 959 611 968 615
rect 794 595 798 599
rect 776 588 780 592
rect 818 588 822 594
rect 776 584 785 588
rect 813 584 822 588
rect 834 589 838 599
rect 873 596 882 600
rect 854 589 858 593
rect 878 590 882 596
rect 895 597 899 601
rect 895 593 905 597
rect 834 585 858 589
rect 776 572 780 584
rect 793 576 805 580
rect 794 565 798 576
rect 818 570 822 584
rect 895 581 899 593
rect 913 585 927 589
rect 951 587 959 603
rect 964 596 968 611
rect 987 614 991 789
rect 1072 770 1076 789
rect 1095 786 1099 789
rect 1119 783 1123 789
rect 1114 779 1123 783
rect 1050 765 1054 769
rect 1050 761 1060 765
rect 1050 749 1054 761
rect 1068 753 1082 757
rect 1106 755 1114 771
rect 1119 764 1123 779
rect 1131 755 1135 789
rect 1162 770 1166 789
rect 1185 786 1189 789
rect 1209 783 1213 789
rect 1204 779 1213 783
rect 1106 751 1135 755
rect 1140 765 1144 769
rect 1140 761 1150 765
rect 1106 749 1114 751
rect 1140 749 1144 761
rect 1158 753 1172 757
rect 1196 755 1204 771
rect 1209 764 1213 779
rect 1253 788 1365 792
rect 1397 788 1455 792
rect 1253 755 1257 788
rect 1338 769 1342 788
rect 1361 785 1365 788
rect 1385 782 1389 788
rect 1380 778 1389 782
rect 1196 751 1257 755
rect 1196 749 1204 751
rect 1090 745 1114 749
rect 1180 745 1204 749
rect 1075 712 1079 737
rect 1106 731 1114 745
rect 1119 723 1123 738
rect 1114 719 1123 723
rect 1095 712 1099 716
rect 1119 713 1123 719
rect 1075 708 1099 712
rect 1165 712 1169 737
rect 1196 731 1204 745
rect 1209 723 1213 738
rect 1204 719 1213 723
rect 1185 712 1189 716
rect 1209 713 1213 719
rect 1165 708 1189 712
rect 1035 700 1059 704
rect 1041 695 1045 700
rect 1049 680 1053 687
rect 1075 680 1079 708
rect 1165 699 1169 708
rect 1165 695 1229 699
rect 1030 676 1034 680
rect 1049 676 1080 680
rect 1049 675 1053 676
rect 1041 662 1045 667
rect 1076 663 1080 676
rect 1037 658 1057 662
rect 1076 659 1103 663
rect 1135 660 1193 663
rect 1076 640 1080 659
rect 1099 656 1103 659
rect 1123 653 1127 659
rect 1118 649 1127 653
rect 1054 635 1058 639
rect 1054 631 1064 635
rect 1054 619 1058 631
rect 1072 623 1086 627
rect 1110 625 1118 641
rect 1123 634 1127 649
rect 1135 625 1139 660
rect 1166 659 1193 660
rect 1166 640 1170 659
rect 1189 656 1193 659
rect 1213 653 1217 659
rect 1208 649 1217 653
rect 1110 621 1139 625
rect 1144 635 1148 639
rect 1144 631 1154 635
rect 1110 619 1118 621
rect 1144 619 1148 631
rect 1162 623 1176 627
rect 1200 625 1208 641
rect 1213 634 1217 649
rect 1225 625 1229 695
rect 1200 621 1229 625
rect 1200 619 1208 621
rect 1094 615 1118 619
rect 1184 615 1208 619
rect 987 610 1044 614
rect 951 583 971 587
rect 951 581 959 583
rect 935 577 959 581
rect 831 571 858 575
rect 831 565 835 571
rect 794 561 835 565
rect 854 568 858 571
rect 878 565 882 571
rect 873 561 882 565
rect 831 552 835 561
rect 809 547 813 551
rect 809 543 819 547
rect 809 531 813 543
rect 827 535 841 539
rect 865 537 873 553
rect 878 546 882 561
rect 920 544 924 569
rect 951 563 959 577
rect 964 555 968 570
rect 959 551 968 555
rect 940 544 944 548
rect 964 545 968 551
rect 920 540 944 544
rect 920 537 924 540
rect 865 533 924 537
rect 987 533 991 610
rect 1017 591 1021 610
rect 1040 607 1044 610
rect 1064 604 1068 610
rect 1059 600 1068 604
rect 995 586 999 590
rect 995 582 1005 586
rect 995 570 999 582
rect 1013 574 1027 578
rect 1051 576 1059 592
rect 1064 585 1068 600
rect 1079 582 1083 607
rect 1110 601 1118 615
rect 1123 593 1127 608
rect 1118 589 1127 593
rect 1099 582 1103 586
rect 1123 583 1127 589
rect 1079 578 1103 582
rect 1169 582 1173 607
rect 1200 601 1208 615
rect 1213 593 1217 608
rect 1208 589 1217 593
rect 1189 582 1193 586
rect 1213 583 1217 589
rect 1169 578 1193 582
rect 1079 576 1083 578
rect 1051 572 1083 576
rect 1051 570 1059 572
rect 1035 566 1059 570
rect 1020 533 1024 558
rect 1051 552 1059 566
rect 1169 569 1173 578
rect 1241 569 1245 751
rect 1169 565 1245 569
rect 1253 613 1257 751
rect 1316 764 1320 768
rect 1316 760 1326 764
rect 1316 748 1320 760
rect 1334 752 1348 756
rect 1372 754 1380 770
rect 1385 763 1389 778
rect 1397 754 1401 788
rect 1428 769 1432 788
rect 1451 785 1455 788
rect 1475 782 1479 788
rect 1470 778 1479 782
rect 1372 750 1401 754
rect 1406 764 1410 768
rect 1406 760 1416 764
rect 1372 748 1380 750
rect 1406 748 1410 760
rect 1424 752 1438 756
rect 1462 754 1470 770
rect 1475 763 1479 778
rect 1462 750 1511 754
rect 1462 748 1470 750
rect 1356 744 1380 748
rect 1446 744 1470 748
rect 1341 711 1345 736
rect 1372 730 1380 744
rect 1385 722 1389 737
rect 1380 718 1389 722
rect 1361 711 1365 715
rect 1385 712 1389 718
rect 1341 707 1365 711
rect 1431 711 1435 736
rect 1462 730 1470 744
rect 1475 722 1479 737
rect 1470 718 1479 722
rect 1451 711 1455 715
rect 1475 712 1479 718
rect 1431 707 1455 711
rect 1341 679 1345 707
rect 1431 698 1435 707
rect 1431 694 1495 698
rect 1337 675 1346 679
rect 1342 662 1346 675
rect 1342 658 1369 662
rect 1401 659 1459 662
rect 1342 639 1346 658
rect 1365 655 1369 658
rect 1389 652 1393 658
rect 1384 648 1393 652
rect 1320 634 1324 638
rect 1320 630 1330 634
rect 1320 618 1324 630
rect 1338 622 1352 626
rect 1376 624 1384 640
rect 1389 633 1393 648
rect 1401 624 1405 659
rect 1432 658 1459 659
rect 1432 639 1436 658
rect 1455 655 1459 658
rect 1479 652 1483 658
rect 1474 648 1483 652
rect 1376 620 1405 624
rect 1410 634 1414 638
rect 1410 630 1420 634
rect 1376 618 1384 620
rect 1410 618 1414 630
rect 1428 622 1442 626
rect 1466 624 1474 640
rect 1479 633 1483 648
rect 1491 624 1495 694
rect 1466 620 1495 624
rect 1466 618 1474 620
rect 1360 614 1384 618
rect 1450 614 1474 618
rect 1253 609 1310 613
rect 1064 544 1068 559
rect 1059 540 1068 544
rect 1040 533 1044 537
rect 1064 534 1068 540
rect 865 531 873 533
rect 849 527 873 531
rect 987 529 1044 533
rect 1253 532 1257 609
rect 1283 590 1287 609
rect 1306 606 1310 609
rect 1330 603 1334 609
rect 1325 599 1334 603
rect 1261 585 1265 589
rect 1261 581 1271 585
rect 1261 569 1265 581
rect 1279 573 1293 577
rect 1317 575 1325 591
rect 1330 584 1334 599
rect 1345 581 1349 606
rect 1376 600 1384 614
rect 1389 592 1393 607
rect 1384 588 1393 592
rect 1365 581 1369 585
rect 1389 582 1393 588
rect 1345 577 1369 581
rect 1435 581 1439 606
rect 1466 600 1474 614
rect 1479 592 1483 607
rect 1474 588 1483 592
rect 1455 581 1459 585
rect 1479 582 1483 588
rect 1435 577 1459 581
rect 1345 575 1349 577
rect 1317 571 1349 575
rect 1317 569 1325 571
rect 1301 565 1325 569
rect 1286 532 1290 557
rect 1317 551 1325 565
rect 1435 568 1439 577
rect 1507 568 1511 750
rect 1435 564 1511 568
rect 1330 543 1334 558
rect 1325 539 1334 543
rect 1306 532 1310 536
rect 1330 533 1334 539
rect 1253 528 1310 532
rect 834 494 838 519
rect 865 513 873 527
rect 878 505 882 520
rect 873 501 882 505
rect 854 494 858 498
rect 878 495 882 501
rect 987 517 1099 521
rect 1131 517 1189 521
rect 764 490 858 494
rect 405 464 461 468
rect 405 462 413 464
rect 389 458 413 462
rect 374 439 378 450
rect 405 444 413 458
rect 457 461 461 464
rect 457 457 484 461
rect 334 435 378 439
rect 418 436 422 451
rect 457 438 461 457
rect 480 454 484 457
rect 504 451 508 457
rect 499 447 508 451
rect 334 431 338 435
rect 316 424 320 428
rect 358 424 362 430
rect 316 420 325 424
rect 353 420 362 424
rect 374 425 378 435
rect 413 432 422 436
rect 394 425 398 429
rect 418 426 422 432
rect 435 433 439 437
rect 435 429 445 433
rect 374 421 398 425
rect 316 408 320 420
rect 333 412 345 416
rect 334 401 338 412
rect 358 406 362 420
rect 435 417 439 429
rect 453 421 467 425
rect 491 423 499 439
rect 504 432 508 447
rect 491 419 514 423
rect 491 417 499 419
rect 475 413 499 417
rect 371 407 398 411
rect 371 401 375 407
rect 334 397 375 401
rect 394 404 398 407
rect 418 401 422 407
rect 413 397 422 401
rect 371 388 375 397
rect 349 383 353 387
rect 349 379 359 383
rect 349 367 353 379
rect 367 371 381 375
rect 405 373 413 389
rect 418 382 422 397
rect 460 380 464 405
rect 491 399 499 413
rect 504 391 508 406
rect 499 387 508 391
rect 480 380 484 384
rect 504 381 508 387
rect 460 376 484 380
rect 460 373 464 376
rect 405 369 464 373
rect 405 367 413 369
rect 389 363 413 367
rect 374 330 378 355
rect 405 349 413 363
rect 418 341 422 356
rect 413 337 422 341
rect 394 330 398 334
rect 418 331 422 337
rect 987 342 991 517
rect 1072 498 1076 517
rect 1095 514 1099 517
rect 1119 511 1123 517
rect 1114 507 1123 511
rect 1050 493 1054 497
rect 1050 489 1060 493
rect 1050 477 1054 489
rect 1068 481 1082 485
rect 1106 483 1114 499
rect 1119 492 1123 507
rect 1131 483 1135 517
rect 1162 498 1166 517
rect 1185 514 1189 517
rect 1209 511 1213 517
rect 1204 507 1213 511
rect 1106 479 1135 483
rect 1140 493 1144 497
rect 1140 489 1150 493
rect 1106 477 1114 479
rect 1140 477 1144 489
rect 1158 481 1172 485
rect 1196 483 1204 499
rect 1209 492 1213 507
rect 1253 516 1365 520
rect 1397 516 1455 520
rect 1253 483 1257 516
rect 1338 497 1342 516
rect 1361 513 1365 516
rect 1385 510 1389 516
rect 1380 506 1389 510
rect 1196 479 1257 483
rect 1196 477 1204 479
rect 1090 473 1114 477
rect 1180 473 1204 477
rect 1075 440 1079 465
rect 1106 459 1114 473
rect 1119 451 1123 466
rect 1114 447 1123 451
rect 1095 440 1099 444
rect 1119 441 1123 447
rect 1075 436 1099 440
rect 1165 440 1169 465
rect 1196 459 1204 473
rect 1209 451 1213 466
rect 1204 447 1213 451
rect 1185 440 1189 444
rect 1209 441 1213 447
rect 1165 436 1189 440
rect 1035 428 1059 432
rect 1041 423 1045 428
rect 1049 408 1053 415
rect 1075 408 1079 436
rect 1165 427 1169 436
rect 1165 423 1229 427
rect 1030 404 1034 408
rect 1049 404 1080 408
rect 1049 403 1053 404
rect 1041 390 1045 395
rect 1076 391 1080 404
rect 1037 386 1057 390
rect 1076 387 1103 391
rect 1135 388 1193 391
rect 1076 368 1080 387
rect 1099 384 1103 387
rect 1123 381 1127 387
rect 1118 377 1127 381
rect 1054 363 1058 367
rect 1054 359 1064 363
rect 1054 347 1058 359
rect 1072 351 1086 355
rect 1110 353 1118 369
rect 1123 362 1127 377
rect 1135 353 1139 388
rect 1166 387 1193 388
rect 1166 368 1170 387
rect 1189 384 1193 387
rect 1213 381 1217 387
rect 1208 377 1217 381
rect 1110 349 1139 353
rect 1144 363 1148 367
rect 1144 359 1154 363
rect 1110 347 1118 349
rect 1144 347 1148 359
rect 1162 351 1176 355
rect 1200 353 1208 369
rect 1213 362 1217 377
rect 1225 353 1229 423
rect 1200 349 1229 353
rect 1200 347 1208 349
rect 1094 343 1118 347
rect 1184 343 1208 347
rect 987 338 1044 342
rect 304 326 398 330
rect 239 306 288 310
rect 239 304 247 306
rect 133 300 157 304
rect 223 300 247 304
rect 118 267 122 292
rect 149 286 157 300
rect 162 278 166 293
rect 157 274 166 278
rect 138 267 142 271
rect 162 268 166 274
rect 118 263 142 267
rect 208 267 212 292
rect 239 286 247 300
rect 252 278 256 293
rect 247 274 256 278
rect 228 267 232 271
rect 252 268 256 274
rect 208 263 232 267
rect 118 235 122 263
rect 208 254 212 263
rect 208 250 272 254
rect 114 231 123 235
rect 119 218 123 231
rect 119 214 146 218
rect 178 215 236 218
rect 119 195 123 214
rect 142 211 146 214
rect 166 208 170 214
rect 161 204 170 208
rect 97 190 101 194
rect 97 186 107 190
rect 97 174 101 186
rect 115 178 129 182
rect 153 180 161 196
rect 166 189 170 204
rect 178 180 182 215
rect 209 214 236 215
rect 209 195 213 214
rect 232 211 236 214
rect 256 208 260 214
rect 251 204 260 208
rect 153 176 182 180
rect 187 190 191 194
rect 187 186 197 190
rect 153 174 161 176
rect 187 174 191 186
rect 205 178 219 182
rect 243 180 251 196
rect 256 189 260 204
rect 268 180 272 250
rect 243 176 272 180
rect 243 174 251 176
rect 137 170 161 174
rect 227 170 251 174
rect 30 165 87 169
rect -159 100 -155 115
rect -164 96 -155 100
rect -183 89 -179 93
rect -159 90 -155 96
rect -236 85 -179 89
rect 30 88 34 165
rect 60 146 64 165
rect 83 162 87 165
rect 107 159 111 165
rect 102 155 111 159
rect 38 141 42 145
rect 38 137 48 141
rect 38 125 42 137
rect 56 129 70 133
rect 94 131 102 147
rect 107 140 111 155
rect 122 137 126 162
rect 153 156 161 170
rect 166 148 170 163
rect 161 144 170 148
rect 142 137 146 141
rect 166 138 170 144
rect 122 133 146 137
rect 212 137 216 162
rect 243 156 251 170
rect 256 148 260 163
rect 251 144 260 148
rect 232 137 236 141
rect 256 138 260 144
rect 212 133 236 137
rect 122 131 126 133
rect 94 127 126 131
rect 94 125 102 127
rect 78 121 102 125
rect 63 88 67 113
rect 94 107 102 121
rect 212 124 216 133
rect 284 124 288 306
rect 326 294 353 298
rect 326 275 330 294
rect 349 291 353 294
rect 373 288 377 294
rect 368 284 377 288
rect 304 270 308 274
rect 304 266 314 270
rect 304 254 308 266
rect 322 258 336 262
rect 360 260 368 276
rect 373 269 377 284
rect 391 280 415 284
rect 397 275 401 280
rect 405 260 409 267
rect 987 261 991 338
rect 1017 319 1021 338
rect 1040 335 1044 338
rect 1064 332 1068 338
rect 1059 328 1068 332
rect 995 314 999 318
rect 995 310 1005 314
rect 995 298 999 310
rect 1013 302 1027 306
rect 1051 304 1059 320
rect 1064 313 1068 328
rect 1079 310 1083 335
rect 1110 329 1118 343
rect 1123 321 1127 336
rect 1118 317 1127 321
rect 1099 310 1103 314
rect 1123 311 1127 317
rect 1079 306 1103 310
rect 1169 310 1173 335
rect 1200 329 1208 343
rect 1213 321 1217 336
rect 1208 317 1217 321
rect 1189 310 1193 314
rect 1213 311 1217 317
rect 1169 306 1193 310
rect 1079 304 1083 306
rect 1051 300 1083 304
rect 1051 298 1059 300
rect 1035 294 1059 298
rect 1020 261 1024 286
rect 1051 280 1059 294
rect 1169 297 1173 306
rect 1241 297 1245 479
rect 1169 293 1245 297
rect 1253 341 1257 479
rect 1316 492 1320 496
rect 1316 488 1326 492
rect 1316 476 1320 488
rect 1334 480 1348 484
rect 1372 482 1380 498
rect 1385 491 1389 506
rect 1397 482 1401 516
rect 1428 497 1432 516
rect 1451 513 1455 516
rect 1475 510 1479 516
rect 1470 506 1479 510
rect 1372 478 1401 482
rect 1406 492 1410 496
rect 1406 488 1416 492
rect 1372 476 1380 478
rect 1406 476 1410 488
rect 1424 480 1438 484
rect 1462 482 1470 498
rect 1475 491 1479 506
rect 1462 478 1511 482
rect 1462 476 1470 478
rect 1356 472 1380 476
rect 1446 472 1470 476
rect 1341 439 1345 464
rect 1372 458 1380 472
rect 1385 450 1389 465
rect 1380 446 1389 450
rect 1361 439 1365 443
rect 1385 440 1389 446
rect 1341 435 1365 439
rect 1431 439 1435 464
rect 1462 458 1470 472
rect 1475 450 1479 465
rect 1470 446 1479 450
rect 1451 439 1455 443
rect 1475 440 1479 446
rect 1431 435 1455 439
rect 1341 407 1345 435
rect 1431 426 1435 435
rect 1431 422 1495 426
rect 1337 403 1346 407
rect 1342 390 1346 403
rect 1342 386 1369 390
rect 1401 387 1459 390
rect 1342 367 1346 386
rect 1365 383 1369 386
rect 1389 380 1393 386
rect 1384 376 1393 380
rect 1320 362 1324 366
rect 1320 358 1330 362
rect 1320 346 1324 358
rect 1338 350 1352 354
rect 1376 352 1384 368
rect 1389 361 1393 376
rect 1401 352 1405 387
rect 1432 386 1459 387
rect 1432 367 1436 386
rect 1455 383 1459 386
rect 1479 380 1483 386
rect 1474 376 1483 380
rect 1376 348 1405 352
rect 1410 362 1414 366
rect 1410 358 1420 362
rect 1376 346 1384 348
rect 1410 346 1414 358
rect 1428 350 1442 354
rect 1466 352 1474 368
rect 1479 361 1483 376
rect 1491 352 1495 422
rect 1466 348 1495 352
rect 1466 346 1474 348
rect 1360 342 1384 346
rect 1450 342 1474 346
rect 1253 337 1310 341
rect 1064 272 1068 287
rect 1059 268 1068 272
rect 1040 261 1044 265
rect 1064 262 1068 268
rect 360 256 390 260
rect 405 256 426 260
rect 987 257 1044 261
rect 1253 260 1257 337
rect 1283 318 1287 337
rect 1306 334 1310 337
rect 1330 331 1334 337
rect 1325 327 1334 331
rect 1261 313 1265 317
rect 1261 309 1271 313
rect 1261 297 1265 309
rect 1279 301 1293 305
rect 1317 303 1325 319
rect 1330 312 1334 327
rect 1345 309 1349 334
rect 1376 328 1384 342
rect 1389 320 1393 335
rect 1384 316 1393 320
rect 1365 309 1369 313
rect 1389 310 1393 316
rect 1345 305 1369 309
rect 1435 309 1439 334
rect 1466 328 1474 342
rect 1479 320 1483 335
rect 1474 316 1483 320
rect 1455 309 1459 313
rect 1479 310 1483 316
rect 1435 305 1459 309
rect 1345 303 1349 305
rect 1317 299 1349 303
rect 1317 297 1325 299
rect 1301 293 1325 297
rect 1286 260 1290 285
rect 1317 279 1325 293
rect 1435 296 1439 305
rect 1507 296 1511 478
rect 1435 292 1511 296
rect 1330 271 1334 286
rect 1325 267 1334 271
rect 1306 260 1310 264
rect 1330 261 1334 267
rect 1253 256 1310 260
rect 360 254 368 256
rect 405 255 409 256
rect 344 250 368 254
rect 329 217 333 242
rect 360 236 368 250
rect 373 228 377 243
rect 397 242 401 247
rect 393 238 413 242
rect 368 224 377 228
rect 349 217 353 221
rect 373 218 377 224
rect 329 213 353 217
rect 212 120 288 124
rect 107 99 111 114
rect 102 95 111 99
rect 83 88 87 92
rect 107 89 111 95
rect 30 84 87 88
rect -236 73 -124 77
rect -92 73 -34 77
rect -236 -102 -232 73
rect -151 54 -147 73
rect -128 70 -124 73
rect -104 67 -100 73
rect -109 63 -100 67
rect -173 49 -169 53
rect -173 45 -163 49
rect -173 33 -169 45
rect -155 37 -141 41
rect -117 39 -109 55
rect -104 48 -100 63
rect -92 39 -88 73
rect -61 54 -57 73
rect -38 70 -34 73
rect -14 67 -10 73
rect -19 63 -10 67
rect -117 35 -88 39
rect -83 49 -79 53
rect -83 45 -73 49
rect -117 33 -109 35
rect -83 33 -79 45
rect -65 37 -51 41
rect -27 39 -19 55
rect -14 48 -10 63
rect 30 72 142 76
rect 174 72 232 76
rect 30 39 34 72
rect 115 53 119 72
rect 138 69 142 72
rect 162 66 166 72
rect 157 62 166 66
rect -27 35 34 39
rect -27 33 -19 35
rect -133 29 -109 33
rect -43 29 -19 33
rect -148 -4 -144 21
rect -117 15 -109 29
rect -104 7 -100 22
rect -109 3 -100 7
rect -128 -4 -124 0
rect -104 -3 -100 3
rect -148 -8 -124 -4
rect -58 -4 -54 21
rect -27 15 -19 29
rect -14 7 -10 22
rect -19 3 -10 7
rect -38 -4 -34 0
rect -14 -3 -10 3
rect -58 -8 -34 -4
rect -188 -16 -164 -12
rect -182 -21 -178 -16
rect -174 -36 -170 -29
rect -148 -36 -144 -8
rect -58 -17 -54 -8
rect -58 -21 6 -17
rect -193 -40 -189 -36
rect -174 -40 -143 -36
rect -174 -41 -170 -40
rect -182 -54 -178 -49
rect -147 -53 -143 -40
rect -186 -58 -166 -54
rect -147 -57 -120 -53
rect -88 -56 -30 -53
rect -147 -76 -143 -57
rect -124 -60 -120 -57
rect -100 -63 -96 -57
rect -105 -67 -96 -63
rect -169 -81 -165 -77
rect -169 -85 -159 -81
rect -169 -97 -165 -85
rect -151 -93 -137 -89
rect -113 -91 -105 -75
rect -100 -82 -96 -67
rect -88 -91 -84 -56
rect -57 -57 -30 -56
rect -57 -76 -53 -57
rect -34 -60 -30 -57
rect -10 -63 -6 -57
rect -15 -67 -6 -63
rect -113 -95 -84 -91
rect -79 -81 -75 -77
rect -79 -85 -69 -81
rect -113 -97 -105 -95
rect -79 -97 -75 -85
rect -61 -93 -47 -89
rect -23 -91 -15 -75
rect -10 -82 -6 -67
rect 2 -91 6 -21
rect -23 -95 6 -91
rect -23 -97 -15 -95
rect -129 -101 -105 -97
rect -39 -101 -15 -97
rect -236 -106 -179 -102
rect -236 -183 -232 -106
rect -206 -125 -202 -106
rect -183 -109 -179 -106
rect -159 -112 -155 -106
rect -164 -116 -155 -112
rect -228 -130 -224 -126
rect -228 -134 -218 -130
rect -228 -146 -224 -134
rect -210 -142 -196 -138
rect -172 -140 -164 -124
rect -159 -131 -155 -116
rect -144 -134 -140 -109
rect -113 -115 -105 -101
rect -100 -123 -96 -108
rect -105 -127 -96 -123
rect -124 -134 -120 -130
rect -100 -133 -96 -127
rect -144 -138 -120 -134
rect -54 -134 -50 -109
rect -23 -115 -15 -101
rect -10 -123 -6 -108
rect -15 -127 -6 -123
rect -34 -134 -30 -130
rect -10 -133 -6 -127
rect -54 -138 -30 -134
rect -144 -140 -140 -138
rect -172 -144 -140 -140
rect -172 -146 -164 -144
rect -188 -150 -164 -146
rect -203 -183 -199 -158
rect -172 -164 -164 -150
rect -54 -147 -50 -138
rect 18 -147 22 35
rect -54 -151 22 -147
rect 30 -103 34 35
rect 93 48 97 52
rect 93 44 103 48
rect 93 32 97 44
rect 111 36 125 40
rect 149 38 157 54
rect 162 47 166 62
rect 174 38 178 72
rect 205 53 209 72
rect 228 69 232 72
rect 252 66 256 72
rect 247 62 256 66
rect 149 34 178 38
rect 183 48 187 52
rect 183 44 193 48
rect 149 32 157 34
rect 183 32 187 44
rect 201 36 215 40
rect 239 38 247 54
rect 252 47 256 62
rect 239 34 288 38
rect 239 32 247 34
rect 133 28 157 32
rect 223 28 247 32
rect 118 -5 122 20
rect 149 14 157 28
rect 162 6 166 21
rect 157 2 166 6
rect 138 -5 142 -1
rect 162 -4 166 2
rect 118 -9 142 -5
rect 208 -5 212 20
rect 239 14 247 28
rect 252 6 256 21
rect 247 2 256 6
rect 228 -5 232 -1
rect 252 -4 256 2
rect 208 -9 232 -5
rect 118 -37 122 -9
rect 208 -18 212 -9
rect 208 -22 272 -18
rect 114 -41 123 -37
rect 119 -54 123 -41
rect 119 -58 146 -54
rect 178 -57 236 -54
rect 119 -77 123 -58
rect 142 -61 146 -58
rect 166 -64 170 -58
rect 161 -68 170 -64
rect 97 -82 101 -78
rect 97 -86 107 -82
rect 97 -98 101 -86
rect 115 -94 129 -90
rect 153 -92 161 -76
rect 166 -83 170 -68
rect 178 -92 182 -57
rect 209 -58 236 -57
rect 209 -77 213 -58
rect 232 -61 236 -58
rect 256 -64 260 -58
rect 251 -68 260 -64
rect 153 -96 182 -92
rect 187 -82 191 -78
rect 187 -86 197 -82
rect 153 -98 161 -96
rect 187 -98 191 -86
rect 205 -94 219 -90
rect 243 -92 251 -76
rect 256 -83 260 -68
rect 268 -92 272 -22
rect 243 -96 272 -92
rect 243 -98 251 -96
rect 137 -102 161 -98
rect 227 -102 251 -98
rect 30 -107 87 -103
rect -159 -172 -155 -157
rect -164 -176 -155 -172
rect -183 -183 -179 -179
rect -159 -182 -155 -176
rect -236 -187 -179 -183
rect 30 -184 34 -107
rect 60 -126 64 -107
rect 83 -110 87 -107
rect 107 -113 111 -107
rect 102 -117 111 -113
rect 38 -131 42 -127
rect 38 -135 48 -131
rect 38 -147 42 -135
rect 56 -143 70 -139
rect 94 -141 102 -125
rect 107 -132 111 -117
rect 122 -135 126 -110
rect 153 -116 161 -102
rect 166 -124 170 -109
rect 161 -128 170 -124
rect 142 -135 146 -131
rect 166 -134 170 -128
rect 122 -139 146 -135
rect 212 -135 216 -110
rect 243 -116 251 -102
rect 256 -124 260 -109
rect 251 -128 260 -124
rect 232 -135 236 -131
rect 256 -134 260 -128
rect 212 -139 236 -135
rect 122 -141 126 -139
rect 94 -145 126 -141
rect 94 -147 102 -145
rect 78 -151 102 -147
rect 63 -184 67 -159
rect 94 -165 102 -151
rect 212 -148 216 -139
rect 284 -148 288 34
rect 212 -152 288 -148
rect 107 -173 111 -158
rect 102 -177 111 -173
rect 83 -184 87 -180
rect 107 -183 111 -177
rect 30 -188 87 -184
<< labels >>
rlabel metal1 351 476 351 476 1 gnd
rlabel metal1 420 434 420 434 7 vdd
rlabel metal1 420 494 420 494 7 vdd
rlabel metal1 351 381 351 381 1 gnd
rlabel metal1 420 339 420 339 7 vdd
rlabel metal1 420 399 420 399 7 vdd
rlabel metal1 506 449 506 449 7 vdd
rlabel metal1 506 389 506 389 7 vdd
rlabel metal1 437 431 437 431 1 gnd
rlabel metal1 306 268 306 268 1 gnd
rlabel metal1 375 226 375 226 7 vdd
rlabel metal1 375 286 375 286 7 vdd
rlabel metal1 399 240 399 240 1 gnd
rlabel metal1 400 282 400 282 1 vdd
rlabel metal1 351 811 351 811 1 gnd
rlabel metal1 420 769 420 769 7 vdd
rlabel metal1 420 829 420 829 7 vdd
rlabel metal1 351 716 351 716 1 gnd
rlabel metal1 420 674 420 674 7 vdd
rlabel metal1 420 734 420 734 7 vdd
rlabel metal1 506 784 506 784 7 vdd
rlabel metal1 506 724 506 724 7 vdd
rlabel metal1 437 766 437 766 1 gnd
rlabel metal1 306 603 306 603 1 gnd
rlabel metal1 375 561 375 561 7 vdd
rlabel metal1 375 621 375 621 7 vdd
rlabel metal1 399 575 399 575 1 gnd
rlabel metal1 400 617 400 617 1 vdd
rlabel metal1 351 1146 351 1146 1 gnd
rlabel metal1 420 1104 420 1104 7 vdd
rlabel metal1 420 1164 420 1164 7 vdd
rlabel metal1 351 1051 351 1051 1 gnd
rlabel metal1 420 1009 420 1009 7 vdd
rlabel metal1 420 1069 420 1069 7 vdd
rlabel metal1 506 1119 506 1119 7 vdd
rlabel metal1 506 1059 506 1059 7 vdd
rlabel metal1 437 1101 437 1101 1 gnd
rlabel metal1 306 938 306 938 1 gnd
rlabel metal1 375 896 375 896 7 vdd
rlabel metal1 375 956 375 956 7 vdd
rlabel metal1 399 910 399 910 1 gnd
rlabel metal1 400 952 400 952 1 vdd
rlabel metal1 400 1287 400 1287 1 vdd
rlabel metal1 399 1245 399 1245 1 gnd
rlabel metal1 375 1291 375 1291 7 vdd
rlabel metal1 375 1231 375 1231 7 vdd
rlabel metal1 306 1273 306 1273 1 gnd
rlabel metal1 437 1436 437 1436 1 gnd
rlabel metal1 506 1394 506 1394 7 vdd
rlabel metal1 506 1454 506 1454 7 vdd
rlabel metal1 420 1404 420 1404 7 vdd
rlabel metal1 420 1344 420 1344 7 vdd
rlabel metal1 351 1386 351 1386 1 gnd
rlabel metal1 420 1499 420 1499 7 vdd
rlabel metal1 420 1439 420 1439 7 vdd
rlabel metal1 351 1481 351 1481 1 gnd
rlabel metal1 328 1301 328 1301 1 ffa0
rlabel metal1 331 1220 331 1220 1 ffb0
rlabel metal1 328 966 328 966 1 ffa1
rlabel metal1 331 885 331 885 1 ffb1
rlabel metal1 328 631 328 631 1 ffa2
rlabel metal1 331 550 331 550 1 ffb2
rlabel metal1 328 296 328 296 1 ffa3
rlabel metal1 331 215 331 215 1 ffb3
rlabel metal1 504 1426 504 1426 1 p0
rlabel metal1 421 1263 421 1263 1 g0
rlabel metal1 504 1091 504 1091 1 p1
rlabel metal1 421 928 421 928 1 g1
rlabel metal1 504 756 504 756 1 p2
rlabel metal1 421 593 421 593 1 g2
rlabel metal1 504 421 504 421 1 p3
rlabel metal1 421 258 421 258 1 g3
rlabel metal1 544 1038 544 1038 5 vdd
rlabel metal1 582 1038 582 1038 5 vdd
rlabel metal1 620 1038 620 1038 5 vdd
rlabel metal1 658 1038 658 1038 5 vdd
rlabel metal1 528 794 528 794 7 gnd
rlabel metal1 515 1014 515 1014 1 clk_mcc
rlabel metal1 527 845 527 845 1 c_in
rlabel metal1 535 874 535 874 1 p0
rlabel metal1 565 885 565 885 1 g0
rlabel metal1 602 896 602 896 1 p1
rlabel metal1 603 926 603 926 1 g1
rlabel metal1 640 937 640 937 1 p2
rlabel metal1 641 967 641 967 1 g2
rlabel metal1 678 978 678 978 1 p3
rlabel metal1 708 979 708 979 1 g3
rlabel metal1 582 895 582 895 1 c1_bar
rlabel metal1 620 936 620 936 1 c2_bar
rlabel metal1 658 977 658 977 1 c3_bar
rlabel metal1 696 1002 696 1002 1 cout_bar
rlabel metal1 727 997 727 997 1 gnd
rlabel metal1 728 1039 728 1039 1 vdd
rlabel metal1 727 940 727 940 1 gnd
rlabel metal1 728 982 728 982 1 vdd
rlabel metal1 727 883 727 883 1 gnd
rlabel metal1 728 925 728 925 1 vdd
rlabel metal1 727 826 727 826 1 gnd
rlabel metal1 728 868 728 868 1 vdd
rlabel metal1 714 1015 714 1015 1 cout_bar
rlabel metal1 746 1015 746 1015 1 cout
rlabel metal1 714 958 714 958 1 c1_bar
rlabel metal1 746 958 746 958 1 c1
rlabel metal1 714 901 714 901 1 c2_bar
rlabel metal1 746 901 746 901 1 c2
rlabel metal1 714 844 714 844 1 c3_bar
rlabel metal1 746 844 746 844 1 c3
rlabel metal1 897 1061 897 1061 1 gnd
rlabel metal1 966 1019 966 1019 7 vdd
rlabel metal1 966 1079 966 1079 7 vdd
rlabel metal1 880 1029 880 1029 7 vdd
rlabel metal1 880 969 880 969 7 vdd
rlabel metal1 811 1011 811 1011 1 gnd
rlabel metal1 880 1124 880 1124 7 vdd
rlabel metal1 880 1064 880 1064 7 vdd
rlabel metal1 811 1106 811 1106 1 gnd
rlabel metal1 897 828 897 828 1 gnd
rlabel metal1 966 786 966 786 7 vdd
rlabel metal1 966 846 966 846 7 vdd
rlabel metal1 880 796 880 796 7 vdd
rlabel metal1 880 736 880 736 7 vdd
rlabel metal1 811 778 811 778 1 gnd
rlabel metal1 880 891 880 891 7 vdd
rlabel metal1 880 831 880 831 7 vdd
rlabel metal1 811 873 811 873 1 gnd
rlabel metal1 811 1339 811 1339 1 gnd
rlabel metal1 880 1297 880 1297 7 vdd
rlabel metal1 880 1357 880 1357 7 vdd
rlabel metal1 811 1244 811 1244 1 gnd
rlabel metal1 880 1202 880 1202 7 vdd
rlabel metal1 880 1262 880 1262 7 vdd
rlabel metal1 966 1312 966 1312 7 vdd
rlabel metal1 966 1252 966 1252 7 vdd
rlabel metal1 897 1294 897 1294 1 gnd
rlabel metal1 897 595 897 595 1 gnd
rlabel metal1 966 553 966 553 7 vdd
rlabel metal1 966 613 966 613 7 vdd
rlabel metal1 880 563 880 563 7 vdd
rlabel metal1 880 503 880 503 7 vdd
rlabel metal1 811 545 811 545 1 gnd
rlabel metal1 880 658 880 658 7 vdd
rlabel metal1 880 598 880 598 7 vdd
rlabel metal1 811 640 811 640 1 gnd
rlabel metal1 360 1426 360 1426 3 vdd
rlabel metal1 318 1427 318 1427 3 gnd
rlabel metal1 318 1092 318 1092 3 gnd
rlabel metal1 360 1091 360 1091 3 vdd
rlabel metal1 360 756 360 756 3 vdd
rlabel metal1 318 757 318 757 3 gnd
rlabel metal1 360 421 360 421 3 vdd
rlabel metal1 318 422 318 422 3 gnd
rlabel metal1 778 1285 778 1285 3 gnd
rlabel metal1 820 1284 820 1284 3 vdd
rlabel metal1 778 1052 778 1052 3 gnd
rlabel metal1 820 1051 820 1051 3 vdd
rlabel metal1 778 819 778 819 3 gnd
rlabel metal1 820 818 820 818 3 vdd
rlabel metal1 778 586 778 586 3 gnd
rlabel metal1 820 585 820 585 3 vdd
rlabel metal1 322 1491 322 1491 1 gnd
rlabel metal1 323 1533 323 1533 1 vdd
rlabel metal1 322 1156 322 1156 1 gnd
rlabel metal1 323 1198 323 1198 1 vdd
rlabel metal1 323 863 323 863 1 vdd
rlabel metal1 322 821 322 821 1 gnd
rlabel metal1 323 528 323 528 1 vdd
rlabel metal1 322 486 322 486 1 gnd
rlabel metal1 783 1391 783 1391 1 vdd
rlabel metal1 782 1349 782 1349 1 gnd
rlabel metal1 782 1116 782 1116 1 gnd
rlabel metal1 783 1158 783 1158 1 vdd
rlabel metal1 782 883 782 883 1 gnd
rlabel metal1 783 925 783 925 1 vdd
rlabel metal1 782 650 782 650 1 gnd
rlabel metal1 783 692 783 692 1 vdd
rlabel metal1 306 1509 306 1509 1 ffa0
rlabel metal1 336 1442 336 1442 1 ffb0
rlabel metal1 306 1174 306 1174 1 ffa1
rlabel metal1 336 1107 336 1107 1 ffb1
rlabel metal1 306 839 306 839 1 ffa2
rlabel metal1 336 772 336 772 1 ffb2
rlabel metal1 306 504 306 504 1 ffa3
rlabel metal1 336 437 336 437 1 ffb3
rlabel metal1 766 1367 766 1367 1 p0
rlabel metal1 796 1300 796 1300 1 cin
rlabel metal1 766 1134 766 1134 1 p1
rlabel metal1 796 1067 796 1067 1 c1
rlabel metal1 766 901 766 901 1 p2
rlabel metal1 796 834 796 834 1 c2
rlabel metal1 766 668 766 668 1 p3
rlabel metal1 796 601 796 601 1 c3
rlabel metal1 966 585 966 585 1 s3
rlabel metal1 966 818 966 818 1 s2
rlabel metal1 966 1051 966 1051 1 s1
rlabel metal1 966 1284 966 1284 1 s0
rlabel metal1 -8 1839 -8 1839 7 vdd
rlabel metal1 -8 1779 -8 1779 7 vdd
rlabel metal1 -77 1821 -77 1821 1 gnd
rlabel metal1 -12 1966 -12 1966 1 vdd
rlabel metal1 -12 1909 -12 1909 1 vdd
rlabel metal1 -81 1947 -81 1947 1 gnd
rlabel metal1 -180 1848 -180 1848 1 gnd
rlabel metal1 -180 1890 -180 1890 1 vdd
rlabel metal1 -167 1821 -167 1821 1 gnd
rlabel metal1 -98 1779 -98 1779 1 vdd
rlabel metal1 -98 1839 -98 1839 1 vdd
rlabel metal1 -102 1915 -102 1915 1 vdd
rlabel metal1 -102 1965 -102 1965 1 vdd
rlabel metal1 -171 1950 -171 1950 1 gnd
rlabel metal1 -157 1790 -157 1790 1 vdd
rlabel metal1 -157 1730 -157 1730 1 vdd
rlabel metal1 -226 1772 -226 1772 1 gnd
rlabel metal1 258 1838 258 1838 7 vdd
rlabel metal1 258 1778 258 1778 7 vdd
rlabel metal1 189 1820 189 1820 1 gnd
rlabel metal1 254 1965 254 1965 1 vdd
rlabel metal1 254 1908 254 1908 1 vdd
rlabel metal1 185 1946 185 1946 1 gnd
rlabel metal1 99 1820 99 1820 1 gnd
rlabel metal1 168 1778 168 1778 1 vdd
rlabel metal1 168 1838 168 1838 1 vdd
rlabel metal1 164 1914 164 1914 1 vdd
rlabel metal1 164 1964 164 1964 1 vdd
rlabel metal1 95 1949 95 1949 1 gnd
rlabel metal1 109 1789 109 1789 1 vdd
rlabel metal1 109 1729 109 1729 1 vdd
rlabel metal1 40 1771 40 1771 1 gnd
rlabel metal1 -8 1567 -8 1567 7 vdd
rlabel metal1 -8 1507 -8 1507 7 vdd
rlabel metal1 -77 1549 -77 1549 1 gnd
rlabel metal1 -12 1694 -12 1694 1 vdd
rlabel metal1 -12 1637 -12 1637 1 vdd
rlabel metal1 -81 1675 -81 1675 1 gnd
rlabel metal1 -180 1576 -180 1576 1 gnd
rlabel metal1 -180 1618 -180 1618 1 vdd
rlabel metal1 -167 1549 -167 1549 1 gnd
rlabel metal1 -98 1507 -98 1507 1 vdd
rlabel metal1 -98 1567 -98 1567 1 vdd
rlabel metal1 -102 1643 -102 1643 1 vdd
rlabel metal1 -102 1693 -102 1693 1 vdd
rlabel metal1 -171 1678 -171 1678 1 gnd
rlabel metal1 -157 1518 -157 1518 1 vdd
rlabel metal1 -157 1458 -157 1458 1 vdd
rlabel metal1 -226 1500 -226 1500 1 gnd
rlabel metal1 258 1566 258 1566 7 vdd
rlabel metal1 258 1506 258 1506 7 vdd
rlabel metal1 189 1548 189 1548 1 gnd
rlabel metal1 254 1693 254 1693 1 vdd
rlabel metal1 254 1636 254 1636 1 vdd
rlabel metal1 185 1674 185 1674 1 gnd
rlabel metal1 99 1548 99 1548 1 gnd
rlabel metal1 168 1506 168 1506 1 vdd
rlabel metal1 168 1566 168 1566 1 vdd
rlabel metal1 164 1642 164 1642 1 vdd
rlabel metal1 164 1692 164 1692 1 vdd
rlabel metal1 95 1677 95 1677 1 gnd
rlabel metal1 109 1517 109 1517 1 vdd
rlabel metal1 109 1457 109 1457 1 vdd
rlabel metal1 40 1499 40 1499 1 gnd
rlabel metal1 -8 1295 -8 1295 7 vdd
rlabel metal1 -8 1235 -8 1235 7 vdd
rlabel metal1 -77 1277 -77 1277 1 gnd
rlabel metal1 -12 1422 -12 1422 1 vdd
rlabel metal1 -12 1365 -12 1365 1 vdd
rlabel metal1 -81 1403 -81 1403 1 gnd
rlabel metal1 -180 1304 -180 1304 1 gnd
rlabel metal1 -180 1346 -180 1346 1 vdd
rlabel metal1 -167 1277 -167 1277 1 gnd
rlabel metal1 -98 1235 -98 1235 1 vdd
rlabel metal1 -98 1295 -98 1295 1 vdd
rlabel metal1 -102 1371 -102 1371 1 vdd
rlabel metal1 -102 1421 -102 1421 1 vdd
rlabel metal1 -171 1406 -171 1406 1 gnd
rlabel metal1 -157 1246 -157 1246 1 vdd
rlabel metal1 -157 1186 -157 1186 1 vdd
rlabel metal1 -226 1228 -226 1228 1 gnd
rlabel metal1 258 1294 258 1294 7 vdd
rlabel metal1 258 1234 258 1234 7 vdd
rlabel metal1 189 1276 189 1276 1 gnd
rlabel metal1 254 1421 254 1421 1 vdd
rlabel metal1 254 1364 254 1364 1 vdd
rlabel metal1 185 1402 185 1402 1 gnd
rlabel metal1 99 1276 99 1276 1 gnd
rlabel metal1 168 1234 168 1234 1 vdd
rlabel metal1 168 1294 168 1294 1 vdd
rlabel metal1 164 1370 164 1370 1 vdd
rlabel metal1 164 1420 164 1420 1 vdd
rlabel metal1 95 1405 95 1405 1 gnd
rlabel metal1 109 1245 109 1245 1 vdd
rlabel metal1 109 1185 109 1185 1 vdd
rlabel metal1 40 1227 40 1227 1 gnd
rlabel metal1 40 955 40 955 1 gnd
rlabel metal1 109 913 109 913 1 vdd
rlabel metal1 109 973 109 973 1 vdd
rlabel metal1 95 1133 95 1133 1 gnd
rlabel metal1 164 1148 164 1148 1 vdd
rlabel metal1 164 1098 164 1098 1 vdd
rlabel metal1 168 1022 168 1022 1 vdd
rlabel metal1 168 962 168 962 1 vdd
rlabel metal1 99 1004 99 1004 1 gnd
rlabel metal1 185 1130 185 1130 1 gnd
rlabel metal1 254 1092 254 1092 1 vdd
rlabel metal1 254 1149 254 1149 1 vdd
rlabel metal1 189 1004 189 1004 1 gnd
rlabel metal1 258 962 258 962 7 vdd
rlabel metal1 258 1022 258 1022 7 vdd
rlabel metal1 -226 956 -226 956 1 gnd
rlabel metal1 -157 914 -157 914 1 vdd
rlabel metal1 -157 974 -157 974 1 vdd
rlabel metal1 -171 1134 -171 1134 1 gnd
rlabel metal1 -102 1149 -102 1149 1 vdd
rlabel metal1 -102 1099 -102 1099 1 vdd
rlabel metal1 -98 1023 -98 1023 1 vdd
rlabel metal1 -98 963 -98 963 1 vdd
rlabel metal1 -167 1005 -167 1005 1 gnd
rlabel metal1 -180 1074 -180 1074 1 vdd
rlabel metal1 -180 1032 -180 1032 1 gnd
rlabel metal1 -81 1131 -81 1131 1 gnd
rlabel metal1 -12 1093 -12 1093 1 vdd
rlabel metal1 -12 1150 -12 1150 1 vdd
rlabel metal1 -77 1005 -77 1005 1 gnd
rlabel metal1 -8 963 -8 963 7 vdd
rlabel metal1 -8 1023 -8 1023 7 vdd
rlabel metal1 -8 751 -8 751 7 vdd
rlabel metal1 -8 691 -8 691 7 vdd
rlabel metal1 -77 733 -77 733 1 gnd
rlabel metal1 -12 878 -12 878 1 vdd
rlabel metal1 -12 821 -12 821 1 vdd
rlabel metal1 -81 859 -81 859 1 gnd
rlabel metal1 -180 760 -180 760 1 gnd
rlabel metal1 -180 802 -180 802 1 vdd
rlabel metal1 -167 733 -167 733 1 gnd
rlabel metal1 -98 691 -98 691 1 vdd
rlabel metal1 -98 751 -98 751 1 vdd
rlabel metal1 -102 827 -102 827 1 vdd
rlabel metal1 -102 877 -102 877 1 vdd
rlabel metal1 -171 862 -171 862 1 gnd
rlabel metal1 -157 702 -157 702 1 vdd
rlabel metal1 -157 642 -157 642 1 vdd
rlabel metal1 -226 684 -226 684 1 gnd
rlabel metal1 258 750 258 750 7 vdd
rlabel metal1 258 690 258 690 7 vdd
rlabel metal1 189 732 189 732 1 gnd
rlabel metal1 254 877 254 877 1 vdd
rlabel metal1 254 820 254 820 1 vdd
rlabel metal1 185 858 185 858 1 gnd
rlabel metal1 99 732 99 732 1 gnd
rlabel metal1 168 690 168 690 1 vdd
rlabel metal1 168 750 168 750 1 vdd
rlabel metal1 164 826 164 826 1 vdd
rlabel metal1 164 876 164 876 1 vdd
rlabel metal1 95 861 95 861 1 gnd
rlabel metal1 109 701 109 701 1 vdd
rlabel metal1 109 641 109 641 1 vdd
rlabel metal1 40 683 40 683 1 gnd
rlabel metal1 -8 479 -8 479 7 vdd
rlabel metal1 -8 419 -8 419 7 vdd
rlabel metal1 -77 461 -77 461 1 gnd
rlabel metal1 -12 606 -12 606 1 vdd
rlabel metal1 -12 549 -12 549 1 vdd
rlabel metal1 -81 587 -81 587 1 gnd
rlabel metal1 -180 488 -180 488 1 gnd
rlabel metal1 -180 530 -180 530 1 vdd
rlabel metal1 -167 461 -167 461 1 gnd
rlabel metal1 -98 419 -98 419 1 vdd
rlabel metal1 -98 479 -98 479 1 vdd
rlabel metal1 -102 555 -102 555 1 vdd
rlabel metal1 -102 605 -102 605 1 vdd
rlabel metal1 -171 590 -171 590 1 gnd
rlabel metal1 -157 430 -157 430 1 vdd
rlabel metal1 -157 370 -157 370 1 vdd
rlabel metal1 -226 412 -226 412 1 gnd
rlabel metal1 258 478 258 478 7 vdd
rlabel metal1 258 418 258 418 7 vdd
rlabel metal1 189 460 189 460 1 gnd
rlabel metal1 254 605 254 605 1 vdd
rlabel metal1 254 548 254 548 1 vdd
rlabel metal1 185 586 185 586 1 gnd
rlabel metal1 99 460 99 460 1 gnd
rlabel metal1 168 418 168 418 1 vdd
rlabel metal1 168 478 168 478 1 vdd
rlabel metal1 164 554 164 554 1 vdd
rlabel metal1 164 604 164 604 1 vdd
rlabel metal1 95 589 95 589 1 gnd
rlabel metal1 109 429 109 429 1 vdd
rlabel metal1 109 369 109 369 1 vdd
rlabel metal1 40 411 40 411 1 gnd
rlabel metal1 -8 207 -8 207 7 vdd
rlabel metal1 -8 147 -8 147 7 vdd
rlabel metal1 -77 189 -77 189 1 gnd
rlabel metal1 -12 334 -12 334 1 vdd
rlabel metal1 -12 277 -12 277 1 vdd
rlabel metal1 -81 315 -81 315 1 gnd
rlabel metal1 -180 216 -180 216 1 gnd
rlabel metal1 -180 258 -180 258 1 vdd
rlabel metal1 -167 189 -167 189 1 gnd
rlabel metal1 -98 147 -98 147 1 vdd
rlabel metal1 -98 207 -98 207 1 vdd
rlabel metal1 -102 283 -102 283 1 vdd
rlabel metal1 -102 333 -102 333 1 vdd
rlabel metal1 -171 318 -171 318 1 gnd
rlabel metal1 -157 158 -157 158 1 vdd
rlabel metal1 -157 98 -157 98 1 vdd
rlabel metal1 -226 140 -226 140 1 gnd
rlabel metal1 258 206 258 206 7 vdd
rlabel metal1 258 146 258 146 7 vdd
rlabel metal1 189 188 189 188 1 gnd
rlabel metal1 254 333 254 333 1 vdd
rlabel metal1 254 276 254 276 1 vdd
rlabel metal1 185 314 185 314 1 gnd
rlabel metal1 99 188 99 188 1 gnd
rlabel metal1 168 146 168 146 1 vdd
rlabel metal1 168 206 168 206 1 vdd
rlabel metal1 164 282 164 282 1 vdd
rlabel metal1 164 332 164 332 1 vdd
rlabel metal1 95 317 95 317 1 gnd
rlabel metal1 109 157 109 157 1 vdd
rlabel metal1 109 97 109 97 1 vdd
rlabel metal1 40 139 40 139 1 gnd
rlabel metal1 40 -133 40 -133 1 gnd
rlabel metal1 109 -175 109 -175 1 vdd
rlabel metal1 109 -115 109 -115 1 vdd
rlabel metal1 95 45 95 45 1 gnd
rlabel metal1 164 60 164 60 1 vdd
rlabel metal1 164 10 164 10 1 vdd
rlabel metal1 168 -66 168 -66 1 vdd
rlabel metal1 168 -126 168 -126 1 vdd
rlabel metal1 99 -84 99 -84 1 gnd
rlabel metal1 185 42 185 42 1 gnd
rlabel metal1 254 4 254 4 1 vdd
rlabel metal1 254 61 254 61 1 vdd
rlabel metal1 189 -84 189 -84 1 gnd
rlabel metal1 258 -126 258 -126 7 vdd
rlabel metal1 258 -66 258 -66 7 vdd
rlabel metal1 -226 -132 -226 -132 1 gnd
rlabel metal1 -157 -174 -157 -174 1 vdd
rlabel metal1 -157 -114 -157 -114 1 vdd
rlabel metal1 -171 46 -171 46 1 gnd
rlabel metal1 -102 61 -102 61 1 vdd
rlabel metal1 -102 11 -102 11 1 vdd
rlabel metal1 -98 -65 -98 -65 1 vdd
rlabel metal1 -98 -125 -98 -125 1 vdd
rlabel metal1 -167 -83 -167 -83 1 gnd
rlabel metal1 -180 -14 -180 -14 1 vdd
rlabel metal1 -180 -56 -180 -56 1 gnd
rlabel metal1 -81 43 -81 43 1 gnd
rlabel metal1 -12 5 -12 5 1 vdd
rlabel metal1 -12 62 -12 62 1 vdd
rlabel metal1 -77 -83 -77 -83 1 gnd
rlabel metal1 -8 -125 -8 -125 7 vdd
rlabel metal1 -8 -65 -8 -65 7 vdd
rlabel metal1 1215 379 1215 379 7 vdd
rlabel metal1 1215 319 1215 319 7 vdd
rlabel metal1 1146 361 1146 361 1 gnd
rlabel metal1 1211 506 1211 506 1 vdd
rlabel metal1 1211 449 1211 449 1 vdd
rlabel metal1 1142 487 1142 487 1 gnd
rlabel metal1 1043 388 1043 388 1 gnd
rlabel metal1 1043 430 1043 430 1 vdd
rlabel metal1 1056 361 1056 361 1 gnd
rlabel metal1 1125 319 1125 319 1 vdd
rlabel metal1 1125 379 1125 379 1 vdd
rlabel metal1 1121 455 1121 455 1 vdd
rlabel metal1 1121 505 1121 505 1 vdd
rlabel metal1 1052 490 1052 490 1 gnd
rlabel metal1 1066 330 1066 330 1 vdd
rlabel metal1 1066 270 1066 270 1 vdd
rlabel metal1 997 312 997 312 1 gnd
rlabel metal1 1481 378 1481 378 7 vdd
rlabel metal1 1481 318 1481 318 7 vdd
rlabel metal1 1412 360 1412 360 1 gnd
rlabel metal1 1477 505 1477 505 1 vdd
rlabel metal1 1477 448 1477 448 1 vdd
rlabel metal1 1408 486 1408 486 1 gnd
rlabel metal1 1322 360 1322 360 1 gnd
rlabel metal1 1391 318 1391 318 1 vdd
rlabel metal1 1391 378 1391 378 1 vdd
rlabel metal1 1387 454 1387 454 1 vdd
rlabel metal1 1387 504 1387 504 1 vdd
rlabel metal1 1318 489 1318 489 1 gnd
rlabel metal1 1332 329 1332 329 1 vdd
rlabel metal1 1332 269 1332 269 1 vdd
rlabel metal1 1263 311 1263 311 1 gnd
rlabel metal1 1263 583 1263 583 1 gnd
rlabel metal1 1332 541 1332 541 1 vdd
rlabel metal1 1332 601 1332 601 1 vdd
rlabel metal1 1318 761 1318 761 1 gnd
rlabel metal1 1387 776 1387 776 1 vdd
rlabel metal1 1387 726 1387 726 1 vdd
rlabel metal1 1391 650 1391 650 1 vdd
rlabel metal1 1391 590 1391 590 1 vdd
rlabel metal1 1322 632 1322 632 1 gnd
rlabel metal1 1408 758 1408 758 1 gnd
rlabel metal1 1477 720 1477 720 1 vdd
rlabel metal1 1477 777 1477 777 1 vdd
rlabel metal1 1412 632 1412 632 1 gnd
rlabel metal1 1481 590 1481 590 7 vdd
rlabel metal1 1481 650 1481 650 7 vdd
rlabel metal1 997 584 997 584 1 gnd
rlabel metal1 1066 542 1066 542 1 vdd
rlabel metal1 1066 602 1066 602 1 vdd
rlabel metal1 1052 762 1052 762 1 gnd
rlabel metal1 1121 777 1121 777 1 vdd
rlabel metal1 1121 727 1121 727 1 vdd
rlabel metal1 1125 651 1125 651 1 vdd
rlabel metal1 1125 591 1125 591 1 vdd
rlabel metal1 1056 633 1056 633 1 gnd
rlabel metal1 1043 702 1043 702 1 vdd
rlabel metal1 1043 660 1043 660 1 gnd
rlabel metal1 1142 759 1142 759 1 gnd
rlabel metal1 1211 721 1211 721 1 vdd
rlabel metal1 1211 778 1211 778 1 vdd
rlabel metal1 1146 633 1146 633 1 gnd
rlabel metal1 1215 591 1215 591 7 vdd
rlabel metal1 1215 651 1215 651 7 vdd
rlabel metal1 1263 855 1263 855 1 gnd
rlabel metal1 1332 813 1332 813 1 vdd
rlabel metal1 1332 873 1332 873 1 vdd
rlabel metal1 1318 1033 1318 1033 1 gnd
rlabel metal1 1387 1048 1387 1048 1 vdd
rlabel metal1 1387 998 1387 998 1 vdd
rlabel metal1 1391 922 1391 922 1 vdd
rlabel metal1 1391 862 1391 862 1 vdd
rlabel metal1 1322 904 1322 904 1 gnd
rlabel metal1 1408 1030 1408 1030 1 gnd
rlabel metal1 1477 992 1477 992 1 vdd
rlabel metal1 1477 1049 1477 1049 1 vdd
rlabel metal1 1412 904 1412 904 1 gnd
rlabel metal1 1481 862 1481 862 7 vdd
rlabel metal1 1481 922 1481 922 7 vdd
rlabel metal1 997 856 997 856 1 gnd
rlabel metal1 1066 814 1066 814 1 vdd
rlabel metal1 1066 874 1066 874 1 vdd
rlabel metal1 1052 1034 1052 1034 1 gnd
rlabel metal1 1121 1049 1121 1049 1 vdd
rlabel metal1 1121 999 1121 999 1 vdd
rlabel metal1 1125 923 1125 923 1 vdd
rlabel metal1 1125 863 1125 863 1 vdd
rlabel metal1 1056 905 1056 905 1 gnd
rlabel metal1 1043 974 1043 974 1 vdd
rlabel metal1 1043 932 1043 932 1 gnd
rlabel metal1 1142 1031 1142 1031 1 gnd
rlabel metal1 1211 993 1211 993 1 vdd
rlabel metal1 1211 1050 1211 1050 1 vdd
rlabel metal1 1146 905 1146 905 1 gnd
rlabel metal1 1215 863 1215 863 7 vdd
rlabel metal1 1215 923 1215 923 7 vdd
rlabel metal1 1263 1127 1263 1127 1 gnd
rlabel metal1 1332 1085 1332 1085 1 vdd
rlabel metal1 1332 1145 1332 1145 1 vdd
rlabel metal1 1318 1305 1318 1305 1 gnd
rlabel metal1 1387 1320 1387 1320 1 vdd
rlabel metal1 1387 1270 1387 1270 1 vdd
rlabel metal1 1391 1194 1391 1194 1 vdd
rlabel metal1 1391 1134 1391 1134 1 vdd
rlabel metal1 1322 1176 1322 1176 1 gnd
rlabel metal1 1408 1302 1408 1302 1 gnd
rlabel metal1 1477 1264 1477 1264 1 vdd
rlabel metal1 1477 1321 1477 1321 1 vdd
rlabel metal1 1412 1176 1412 1176 1 gnd
rlabel metal1 1481 1134 1481 1134 7 vdd
rlabel metal1 1481 1194 1481 1194 7 vdd
rlabel metal1 997 1128 997 1128 1 gnd
rlabel metal1 1066 1086 1066 1086 1 vdd
rlabel metal1 1066 1146 1066 1146 1 vdd
rlabel metal1 1052 1306 1052 1306 1 gnd
rlabel metal1 1121 1321 1121 1321 1 vdd
rlabel metal1 1121 1271 1121 1271 1 vdd
rlabel metal1 1125 1195 1125 1195 1 vdd
rlabel metal1 1125 1135 1125 1135 1 vdd
rlabel metal1 1056 1177 1056 1177 1 gnd
rlabel metal1 1043 1246 1043 1246 1 vdd
rlabel metal1 1043 1204 1043 1204 1 gnd
rlabel metal1 1142 1303 1142 1303 1 gnd
rlabel metal1 1211 1265 1211 1265 1 vdd
rlabel metal1 1211 1322 1211 1322 1 vdd
rlabel metal1 1146 1177 1146 1177 1 gnd
rlabel metal1 1215 1135 1215 1135 7 vdd
rlabel metal1 1215 1195 1215 1195 7 vdd
rlabel metal1 1215 1467 1215 1467 7 vdd
rlabel metal1 1215 1407 1215 1407 7 vdd
rlabel metal1 1146 1449 1146 1449 1 gnd
rlabel metal1 1211 1594 1211 1594 1 vdd
rlabel metal1 1211 1537 1211 1537 1 vdd
rlabel metal1 1142 1575 1142 1575 1 gnd
rlabel metal1 1043 1476 1043 1476 1 gnd
rlabel metal1 1043 1518 1043 1518 1 vdd
rlabel metal1 1056 1449 1056 1449 1 gnd
rlabel metal1 1125 1407 1125 1407 1 vdd
rlabel metal1 1125 1467 1125 1467 1 vdd
rlabel metal1 1121 1543 1121 1543 1 vdd
rlabel metal1 1121 1593 1121 1593 1 vdd
rlabel metal1 1052 1578 1052 1578 1 gnd
rlabel metal1 1066 1418 1066 1418 1 vdd
rlabel metal1 1066 1358 1066 1358 1 vdd
rlabel metal1 997 1400 997 1400 1 gnd
rlabel metal1 1481 1466 1481 1466 7 vdd
rlabel metal1 1481 1406 1481 1406 7 vdd
rlabel metal1 1412 1448 1412 1448 1 gnd
rlabel metal1 1477 1593 1477 1593 1 vdd
rlabel metal1 1477 1536 1477 1536 1 vdd
rlabel metal1 1408 1574 1408 1574 1 gnd
rlabel metal1 1322 1448 1322 1448 1 gnd
rlabel metal1 1391 1406 1391 1406 1 vdd
rlabel metal1 1391 1466 1391 1466 1 vdd
rlabel metal1 1387 1542 1387 1542 1 vdd
rlabel metal1 1387 1592 1387 1592 1 vdd
rlabel metal1 1318 1577 1318 1577 1 gnd
rlabel metal1 1332 1417 1332 1417 1 vdd
rlabel metal1 1332 1357 1332 1357 1 vdd
rlabel metal1 1263 1399 1263 1399 1 gnd
rlabel metal1 -191 1866 -191 1866 1 clk
rlabel metal1 -191 1594 -191 1594 1 clk
rlabel metal1 -191 1322 -191 1322 1 clk
rlabel metal1 -191 1050 -191 1050 1 clk
rlabel metal1 -191 778 -191 778 1 clk
rlabel metal1 -191 506 -191 506 1 clk
rlabel metal1 -191 234 -191 234 1 clk
rlabel metal1 -191 -38 -191 -38 1 clk
rlabel metal1 116 1865 116 1865 1 clk
rlabel metal1 116 1593 116 1593 1 clk
rlabel metal1 116 1321 116 1321 1 clk
rlabel metal1 116 1049 116 1049 1 clk
rlabel metal1 116 777 116 777 1 clk
rlabel metal1 116 505 116 505 1 clk
rlabel metal1 116 233 116 233 1 clk
rlabel metal1 116 -39 116 -39 1 clk
rlabel metal1 1032 1494 1032 1494 1 clk
rlabel metal1 1032 1222 1032 1222 1 clk
rlabel metal1 1032 950 1032 950 1 clk
rlabel metal1 1032 678 1032 678 1 clk
rlabel metal1 1032 406 1032 406 1 clk
rlabel metal1 1339 405 1339 405 1 clk
rlabel metal1 1339 677 1339 677 1 clk
rlabel metal1 1339 949 1339 949 1 clk
rlabel metal1 1339 1221 1339 1221 1 clk
rlabel metal1 1339 1493 1339 1493 1 clk
rlabel metal1 -234 1979 -234 1979 4 a0
rlabel metal1 -234 1707 -234 1707 3 a1
rlabel metal1 -234 1435 -234 1435 3 a2
rlabel metal1 -234 1163 -234 1163 3 a3
rlabel metal1 -234 891 -234 891 3 b0
rlabel metal1 -234 619 -234 619 3 b1
rlabel metal1 -234 347 -234 347 3 b2
rlabel metal1 -234 75 -234 75 3 b3
rlabel metal1 286 1940 286 1940 1 ffa0
rlabel metal1 270 1810 270 1810 1 ffa0_bar
rlabel metal1 286 1668 286 1668 1 ffa1
rlabel metal1 270 1538 270 1538 1 ffa1_bar
rlabel metal1 286 1396 286 1396 1 ffa2
rlabel metal1 270 1266 270 1266 1 ffa2_bar
rlabel metal1 286 1124 286 1124 1 ffa3
rlabel metal1 270 994 270 994 1 ffa3_bar
rlabel metal1 286 852 286 852 1 ffb0
rlabel metal1 270 722 270 722 1 ffb0_bar
rlabel metal1 286 580 286 580 1 ffb1
rlabel metal1 270 450 270 450 1 ffb1_bar
rlabel metal1 286 308 286 308 1 ffb2
rlabel metal1 270 178 270 178 1 ffb2_bar
rlabel metal1 286 36 286 36 1 ffb3
rlabel metal1 270 -94 270 -94 1 ffb3_bar
rlabel metal1 989 1607 989 1607 1 cout
rlabel metal1 989 1335 989 1335 1 s0
rlabel metal1 989 1063 989 1063 1 s1
rlabel metal1 989 791 989 791 1 s2
rlabel metal1 989 519 989 519 1 s3
rlabel metal1 1509 1568 1509 1568 7 ffcout
rlabel metal1 1493 1438 1493 1438 1 ffcout_bar
rlabel metal1 1509 1296 1509 1296 7 ffs0
rlabel metal1 1493 1166 1493 1166 1 ffs0_bar
rlabel metal1 1509 1024 1509 1024 7 ffs1
rlabel metal1 1493 894 1493 894 1 ffs1_bar
rlabel metal1 1509 752 1509 752 7 ffs2
rlabel metal1 1493 622 1493 622 1 ffs2_bar
rlabel metal1 1509 480 1509 480 7 ffs3
rlabel metal1 1493 350 1493 350 1 ffs3_bar
<< end >>
